-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08087fe",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"97a87383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02f4050d",
    30 => x"74767181",
    31 => x"ff06c80c",
    32 => x"535383ff",
    33 => x"f09c0885",
    34 => x"3871892b",
    35 => x"5271982a",
    36 => x"c80c7190",
    37 => x"2a7081ff",
    38 => x"06c80c51",
    39 => x"71882a70",
    40 => x"81ff06c8",
    41 => x"0c517181",
    42 => x"ff06c80c",
    43 => x"72902a70",
    44 => x"81ff06c8",
    45 => x"0c51c808",
    46 => x"7081ff06",
    47 => x"515182b8",
    48 => x"bf527081",
    49 => x"ff2e0981",
    50 => x"06943881",
    51 => x"ff0bc80c",
    52 => x"c8087081",
    53 => x"ff06ff14",
    54 => x"54515171",
    55 => x"e5387083",
    56 => x"ffe0800c",
    57 => x"028c050d",
    58 => x"0402fc05",
    59 => x"0d81c751",
    60 => x"81ff0bc8",
    61 => x"0cff1151",
    62 => x"708025f4",
    63 => x"38028405",
    64 => x"0d0402f0",
    65 => x"050da080",
    66 => x"81e92d81",
    67 => x"9c9f5380",
    68 => x"5287fc80",
    69 => x"f751a080",
    70 => x"80f42d83",
    71 => x"ffe08008",
    72 => x"5483ffe0",
    73 => x"8008812e",
    74 => x"098106ab",
    75 => x"3881ff0b",
    76 => x"c80c820a",
    77 => x"52849c80",
    78 => x"e951a080",
    79 => x"80f42d83",
    80 => x"ffe08008",
    81 => x"8d3881ff",
    82 => x"0bc80c73",
    83 => x"53a08082",
    84 => x"de04a080",
    85 => x"81e92dff",
    86 => x"135372ff",
    87 => x"b2387283",
    88 => x"ffe0800c",
    89 => x"0290050d",
    90 => x"0402f405",
    91 => x"0d81ff0b",
    92 => x"c80c9353",
    93 => x"805287fc",
    94 => x"80c151a0",
    95 => x"8080f42d",
    96 => x"83ffe080",
    97 => x"088d3881",
    98 => x"ff0bc80c",
    99 => x"8153a080",
   100 => x"839e04a0",
   101 => x"8081e92d",
   102 => x"ff135372",
   103 => x"d7387283",
   104 => x"ffe0800c",
   105 => x"028c050d",
   106 => x"0402f005",
   107 => x"0da08081",
   108 => x"e92d83aa",
   109 => x"52849c80",
   110 => x"c851a080",
   111 => x"80f42d83",
   112 => x"ffe08008",
   113 => x"812e0981",
   114 => x"069038cc",
   115 => x"087083ff",
   116 => x"ff065153",
   117 => x"7283aa2e",
   118 => x"9938a080",
   119 => x"82e92da0",
   120 => x"8083eb04",
   121 => x"8154a080",
   122 => x"84cc0480",
   123 => x"54a08084",
   124 => x"cc0481ff",
   125 => x"0bc80cb1",
   126 => x"53a08082",
   127 => x"822d83ff",
   128 => x"e0800880",
   129 => x"2eb73880",
   130 => x"5287fc80",
   131 => x"fa51a080",
   132 => x"80f42d83",
   133 => x"ffe08008",
   134 => x"a43881ff",
   135 => x"0bc80cc8",
   136 => x"08cc0871",
   137 => x"862a7081",
   138 => x"0683ffe0",
   139 => x"80085351",
   140 => x"52555372",
   141 => x"802e9538",
   142 => x"a08083e4",
   143 => x"0472822e",
   144 => x"ffa938ff",
   145 => x"135372ff",
   146 => x"b0387254",
   147 => x"7383ffe0",
   148 => x"800c0290",
   149 => x"050d0402",
   150 => x"f4050d81",
   151 => x"0b83fff0",
   152 => x"9c0cc408",
   153 => x"708f2a70",
   154 => x"81065151",
   155 => x"5372f338",
   156 => x"72c40ca0",
   157 => x"8081e92d",
   158 => x"c408708f",
   159 => x"2a708106",
   160 => x"51515372",
   161 => x"f338810b",
   162 => x"c40c8753",
   163 => x"805284d4",
   164 => x"80c051a0",
   165 => x"8080f42d",
   166 => x"83ffe080",
   167 => x"08812e96",
   168 => x"3872822e",
   169 => x"09810688",
   170 => x"388053a0",
   171 => x"8085ee04",
   172 => x"ff135372",
   173 => x"d738a080",
   174 => x"83a92d83",
   175 => x"ffe08008",
   176 => x"83fff09c",
   177 => x"0c815287",
   178 => x"fc80d051",
   179 => x"a08080f4",
   180 => x"2d81ff0b",
   181 => x"c80cc408",
   182 => x"708f2a70",
   183 => x"81065151",
   184 => x"5372f338",
   185 => x"72c40c81",
   186 => x"ff0bc80c",
   187 => x"81537283",
   188 => x"ffe0800c",
   189 => x"028c050d",
   190 => x"04800b83",
   191 => x"ffe0800c",
   192 => x"0402e805",
   193 => x"0d785580",
   194 => x"56c40870",
   195 => x"8f2a7081",
   196 => x"06515153",
   197 => x"72f33882",
   198 => x"810bc40c",
   199 => x"81ff0bc8",
   200 => x"0c775287",
   201 => x"fc80d151",
   202 => x"a08080f4",
   203 => x"2d83ffe0",
   204 => x"800880d2",
   205 => x"3880dbc6",
   206 => x"df5481ff",
   207 => x"0bc80cc8",
   208 => x"087081ff",
   209 => x"06515372",
   210 => x"81fe2e09",
   211 => x"81069b38",
   212 => x"80ff54cc",
   213 => x"08757084",
   214 => x"05570cff",
   215 => x"14547380",
   216 => x"25f13881",
   217 => x"56a08086",
   218 => x"f004ff14",
   219 => x"5473cb38",
   220 => x"81ff0bc8",
   221 => x"0cc40870",
   222 => x"8f2a7081",
   223 => x"06515153",
   224 => x"72f33872",
   225 => x"c40c7583",
   226 => x"ffe0800c",
   227 => x"0298050d",
   228 => x"0402f405",
   229 => x"0d747088",
   230 => x"2a83fe80",
   231 => x"06707298",
   232 => x"2a077288",
   233 => x"2b87fc80",
   234 => x"80067398",
   235 => x"2b81f00a",
   236 => x"06717307",
   237 => x"0783ffe0",
   238 => x"800c5651",
   239 => x"5351028c",
   240 => x"050d0402",
   241 => x"f4050d02",
   242 => x"9205a080",
   243 => x"809f2d70",
   244 => x"882a7188",
   245 => x"2b077083",
   246 => x"ffff0683",
   247 => x"ffe0800c",
   248 => x"5252028c",
   249 => x"050d0402",
   250 => x"f8050d73",
   251 => x"70902b71",
   252 => x"902a0783",
   253 => x"ffe0800c",
   254 => x"52028805",
   255 => x"0d0402ec",
   256 => x"050d88bd",
   257 => x"0bff880c",
   258 => x"800b870a",
   259 => x"0cf80883",
   260 => x"fff0900c",
   261 => x"fc0883ff",
   262 => x"f0940c84",
   263 => x"eacda880",
   264 => x"0b83fff0",
   265 => x"980ca080",
   266 => x"84d72d83",
   267 => x"ffe08008",
   268 => x"902b7090",
   269 => x"2c515372",
   270 => x"802e81d1",
   271 => x"38a0808a",
   272 => x"e12d83ff",
   273 => x"e0905283",
   274 => x"fff09051",
   275 => x"a08095f2",
   276 => x"2d83ffe0",
   277 => x"8008802e",
   278 => x"81b33883",
   279 => x"ffe09054",
   280 => x"80557370",
   281 => x"810555a0",
   282 => x"8080b42d",
   283 => x"5372a02e",
   284 => x"80de3872",
   285 => x"a32e80fd",
   286 => x"387280c7",
   287 => x"2e098106",
   288 => x"8b38a080",
   289 => x"80882da0",
   290 => x"8089ac04",
   291 => x"728a2e09",
   292 => x"81068b38",
   293 => x"a0808090",
   294 => x"2da08089",
   295 => x"ac047280",
   296 => x"cc2e0981",
   297 => x"06863883",
   298 => x"ffe09054",
   299 => x"7281df06",
   300 => x"f0057081",
   301 => x"ff065153",
   302 => x"b8732789",
   303 => x"38ef1370",
   304 => x"81ff0651",
   305 => x"5374842b",
   306 => x"730755a0",
   307 => x"8088e204",
   308 => x"72a32ea1",
   309 => x"38737081",
   310 => x"0555a080",
   311 => x"80b42d53",
   312 => x"72a02ef1",
   313 => x"38ff1475",
   314 => x"53705254",
   315 => x"a08095f2",
   316 => x"2d74870a",
   317 => x"0c737081",
   318 => x"0555a080",
   319 => x"80b42d53",
   320 => x"728a2e09",
   321 => x"8106ee38",
   322 => x"a08088e0",
   323 => x"04800b83",
   324 => x"ffe0800c",
   325 => x"0294050d",
   326 => x"0402e805",
   327 => x"0d77797b",
   328 => x"58555580",
   329 => x"53727625",
   330 => x"ab387470",
   331 => x"810556a0",
   332 => x"8080b42d",
   333 => x"74708105",
   334 => x"56a08080",
   335 => x"b42d5252",
   336 => x"71712e88",
   337 => x"388151a0",
   338 => x"808ad604",
   339 => x"811353a0",
   340 => x"808aa504",
   341 => x"80517083",
   342 => x"ffe0800c",
   343 => x"0298050d",
   344 => x"0402d805",
   345 => x"0dff0b83",
   346 => x"fff4c80c",
   347 => x"800b83ff",
   348 => x"f4dc0c83",
   349 => x"fff0b452",
   350 => x"8051a080",
   351 => x"86812d83",
   352 => x"ffe08008",
   353 => x"902b7090",
   354 => x"2c705751",
   355 => x"5473802e",
   356 => x"86d73880",
   357 => x"56810b83",
   358 => x"fff0a80c",
   359 => x"8853a080",
   360 => x"97b85283",
   361 => x"fff0ea51",
   362 => x"a0808a99",
   363 => x"2d83ffe0",
   364 => x"8008762e",
   365 => x"0981068b",
   366 => x"3883ffe0",
   367 => x"800883ff",
   368 => x"f0a80c88",
   369 => x"53a08097",
   370 => x"c45283ff",
   371 => x"f18651a0",
   372 => x"808a992d",
   373 => x"83ffe080",
   374 => x"088b3883",
   375 => x"ffe08008",
   376 => x"83fff0a8",
   377 => x"0c83fff0",
   378 => x"a808802e",
   379 => x"81a03883",
   380 => x"fff3fa0b",
   381 => x"a08080b4",
   382 => x"2d83fff3",
   383 => x"fb0ba080",
   384 => x"80b42d71",
   385 => x"982b7190",
   386 => x"2b0783ff",
   387 => x"f3fc0ba0",
   388 => x"8080b42d",
   389 => x"70882b72",
   390 => x"0783fff3",
   391 => x"fd0ba080",
   392 => x"80b42d71",
   393 => x"0783fff4",
   394 => x"b20ba080",
   395 => x"80b42d83",
   396 => x"fff4b30b",
   397 => x"a08080b4",
   398 => x"2d71882b",
   399 => x"07535f54",
   400 => x"525a5657",
   401 => x"557381ab",
   402 => x"aa2e0981",
   403 => x"06933875",
   404 => x"51a08087",
   405 => x"912d83ff",
   406 => x"e0800856",
   407 => x"a0808cee",
   408 => x"04805573",
   409 => x"82d4d52e",
   410 => x"09810684",
   411 => x"fc3883ff",
   412 => x"f0b45275",
   413 => x"51a08086",
   414 => x"812d83ff",
   415 => x"e0800890",
   416 => x"2b70902c",
   417 => x"70575154",
   418 => x"73802e84",
   419 => x"dc388853",
   420 => x"a08097c4",
   421 => x"5283fff1",
   422 => x"8651a080",
   423 => x"8a992d83",
   424 => x"ffe08008",
   425 => x"8d38810b",
   426 => x"83fff4dc",
   427 => x"0ca0808d",
   428 => x"d2048853",
   429 => x"a08097b8",
   430 => x"5283fff0",
   431 => x"ea51a080",
   432 => x"8a992d80",
   433 => x"5583ffe0",
   434 => x"8008752e",
   435 => x"09810684",
   436 => x"983883ff",
   437 => x"f4b20ba0",
   438 => x"8080b42d",
   439 => x"547380d5",
   440 => x"2e098106",
   441 => x"80db3883",
   442 => x"fff4b30b",
   443 => x"a08080b4",
   444 => x"2d547381",
   445 => x"aa2e0981",
   446 => x"0680c638",
   447 => x"800b83ff",
   448 => x"f0b40ba0",
   449 => x"8080b42d",
   450 => x"56547481",
   451 => x"e92e8338",
   452 => x"81547481",
   453 => x"eb2e8c38",
   454 => x"80557375",
   455 => x"2e098106",
   456 => x"83c73883",
   457 => x"fff0bf0b",
   458 => x"a08080b4",
   459 => x"2d557491",
   460 => x"3883fff0",
   461 => x"c00ba080",
   462 => x"80b42d54",
   463 => x"73822e88",
   464 => x"388055a0",
   465 => x"8091e904",
   466 => x"83fff0c1",
   467 => x"0ba08080",
   468 => x"b42d7083",
   469 => x"fff4e40c",
   470 => x"ff0583ff",
   471 => x"f4d80c83",
   472 => x"fff0c20b",
   473 => x"a08080b4",
   474 => x"2d83fff0",
   475 => x"c30ba080",
   476 => x"80b42d58",
   477 => x"76057782",
   478 => x"80290570",
   479 => x"83fff4cc",
   480 => x"0c83fff0",
   481 => x"c40ba080",
   482 => x"80b42d70",
   483 => x"83fff4c4",
   484 => x"0c83fff4",
   485 => x"dc085957",
   486 => x"5876802e",
   487 => x"81df3888",
   488 => x"53a08097",
   489 => x"c45283ff",
   490 => x"f18651a0",
   491 => x"808a992d",
   492 => x"83ffe080",
   493 => x"0882b238",
   494 => x"83fff4e4",
   495 => x"0870842b",
   496 => x"83fff4b4",
   497 => x"0c7083ff",
   498 => x"f4e00c83",
   499 => x"fff0d90b",
   500 => x"a08080b4",
   501 => x"2d83fff0",
   502 => x"d80ba080",
   503 => x"80b42d71",
   504 => x"82802905",
   505 => x"83fff0da",
   506 => x"0ba08080",
   507 => x"b42d7084",
   508 => x"80802912",
   509 => x"83fff0db",
   510 => x"0ba08080",
   511 => x"b42d7081",
   512 => x"800a2912",
   513 => x"7083fff0",
   514 => x"ac0c83ff",
   515 => x"f4c40871",
   516 => x"2983fff4",
   517 => x"cc080570",
   518 => x"83fff4ec",
   519 => x"0c83fff0",
   520 => x"e10ba080",
   521 => x"80b42d83",
   522 => x"fff0e00b",
   523 => x"a08080b4",
   524 => x"2d718280",
   525 => x"290583ff",
   526 => x"f0e20ba0",
   527 => x"8080b42d",
   528 => x"70848080",
   529 => x"291283ff",
   530 => x"f0e30ba0",
   531 => x"8080b42d",
   532 => x"70982b81",
   533 => x"f00a0672",
   534 => x"057083ff",
   535 => x"f0b00cfe",
   536 => x"117e2977",
   537 => x"0583fff4",
   538 => x"d40c5259",
   539 => x"5243545e",
   540 => x"51525952",
   541 => x"5d575957",
   542 => x"a08091e7",
   543 => x"0483fff0",
   544 => x"c60ba080",
   545 => x"80b42d83",
   546 => x"fff0c50b",
   547 => x"a08080b4",
   548 => x"2d718280",
   549 => x"29057083",
   550 => x"fff4b40c",
   551 => x"70a02983",
   552 => x"ff057089",
   553 => x"2a7083ff",
   554 => x"f4e00c83",
   555 => x"fff0cb0b",
   556 => x"a08080b4",
   557 => x"2d83fff0",
   558 => x"ca0ba080",
   559 => x"80b42d71",
   560 => x"82802905",
   561 => x"7083fff0",
   562 => x"ac0c7b71",
   563 => x"291e7083",
   564 => x"fff4d40c",
   565 => x"7d83fff0",
   566 => x"b00c7305",
   567 => x"83fff4ec",
   568 => x"0c555e51",
   569 => x"51555581",
   570 => x"557483ff",
   571 => x"e0800c02",
   572 => x"a8050d04",
   573 => x"02e8050d",
   574 => x"7770872c",
   575 => x"7180ff06",
   576 => x"56565383",
   577 => x"fff4dc08",
   578 => x"8a387288",
   579 => x"2c7381ff",
   580 => x"06555574",
   581 => x"83fff4c8",
   582 => x"082eac38",
   583 => x"83fff0b4",
   584 => x"5283fff4",
   585 => x"cc081551",
   586 => x"a0808681",
   587 => x"2d83ffe0",
   588 => x"8008902b",
   589 => x"70902c70",
   590 => x"58515372",
   591 => x"802e80cb",
   592 => x"387483ff",
   593 => x"f4c80c83",
   594 => x"fff4dc08",
   595 => x"802ea038",
   596 => x"73842983",
   597 => x"fff0b405",
   598 => x"70085253",
   599 => x"a0808791",
   600 => x"2d83ffe0",
   601 => x"8008f00a",
   602 => x"0654a080",
   603 => x"93890473",
   604 => x"1083fff0",
   605 => x"b40570a0",
   606 => x"80809f2d",
   607 => x"5253a080",
   608 => x"87c32d83",
   609 => x"ffe08008",
   610 => x"54735675",
   611 => x"83ffe080",
   612 => x"0c029805",
   613 => x"0d0402cc",
   614 => x"050d7e60",
   615 => x"5e5b8056",
   616 => x"ff0b83ff",
   617 => x"f4c80c83",
   618 => x"fff0b008",
   619 => x"83fff4d4",
   620 => x"08565a83",
   621 => x"fff4dc08",
   622 => x"762e8e38",
   623 => x"83fff4e4",
   624 => x"08842b58",
   625 => x"a08093d1",
   626 => x"0483fff4",
   627 => x"e008842b",
   628 => x"58805978",
   629 => x"782781c9",
   630 => x"38788f06",
   631 => x"a0175754",
   632 => x"73953883",
   633 => x"fff0b452",
   634 => x"74518115",
   635 => x"55a08086",
   636 => x"812d83ff",
   637 => x"f0b45680",
   638 => x"76a08080",
   639 => x"b42d5557",
   640 => x"73772e83",
   641 => x"38815773",
   642 => x"81e52e81",
   643 => x"8c388170",
   644 => x"7806555c",
   645 => x"73802e81",
   646 => x"80388b16",
   647 => x"a08080b4",
   648 => x"2d980657",
   649 => x"7680f238",
   650 => x"8b537c52",
   651 => x"7551a080",
   652 => x"8a992d83",
   653 => x"ffe08008",
   654 => x"80df389c",
   655 => x"160851a0",
   656 => x"8087912d",
   657 => x"83ffe080",
   658 => x"08841c0c",
   659 => x"9a16a080",
   660 => x"809f2d51",
   661 => x"a08087c3",
   662 => x"2d83ffe0",
   663 => x"800883ff",
   664 => x"e0800855",
   665 => x"5583fff4",
   666 => x"dc08802e",
   667 => x"9e389416",
   668 => x"a080809f",
   669 => x"2d51a080",
   670 => x"87c32d83",
   671 => x"ffe08008",
   672 => x"902b83ff",
   673 => x"f00a0670",
   674 => x"16515473",
   675 => x"881c0c76",
   676 => x"7b0c7b54",
   677 => x"a08095e7",
   678 => x"04811959",
   679 => x"a08093d3",
   680 => x"0483fff4",
   681 => x"dc08802e",
   682 => x"bc387951",
   683 => x"a08091f4",
   684 => x"2d83ffe0",
   685 => x"800883ff",
   686 => x"e0800880",
   687 => x"fffffff8",
   688 => x"06555a73",
   689 => x"80ffffff",
   690 => x"f82e9a38",
   691 => x"83ffe080",
   692 => x"08fe0583",
   693 => x"fff4e408",
   694 => x"2983fff4",
   695 => x"ec080555",
   696 => x"a08093d1",
   697 => x"04805473",
   698 => x"83ffe080",
   699 => x"0c02b405",
   700 => x"0d0402e4",
   701 => x"050d7979",
   702 => x"5383fff4",
   703 => x"b85255a0",
   704 => x"8093962d",
   705 => x"83ffe080",
   706 => x"0881ff06",
   707 => x"70555372",
   708 => x"802e8189",
   709 => x"3883fff4",
   710 => x"bc0883ff",
   711 => x"05892a57",
   712 => x"80705556",
   713 => x"75772580",
   714 => x"f23883ff",
   715 => x"f4c008fe",
   716 => x"0583fff4",
   717 => x"e4082983",
   718 => x"fff4ec08",
   719 => x"117583ff",
   720 => x"f4d80806",
   721 => x"05765452",
   722 => x"53a08086",
   723 => x"812d83ff",
   724 => x"e0800890",
   725 => x"2b70902c",
   726 => x"51537280",
   727 => x"2eb63881",
   728 => x"147083ff",
   729 => x"f4d80806",
   730 => x"54547296",
   731 => x"3883fff4",
   732 => x"c00851a0",
   733 => x"8091f42d",
   734 => x"83ffe080",
   735 => x"0883fff4",
   736 => x"c00c8480",
   737 => x"15811757",
   738 => x"55767624",
   739 => x"ff9c38a0",
   740 => x"80979b04",
   741 => x"7254a080",
   742 => x"979d0481",
   743 => x"547383ff",
   744 => x"e0800c02",
   745 => x"9c050d04",
   746 => x"00ffffff",
   747 => x"ff00ffff",
   748 => x"ffff00ff",
   749 => x"ffffff00",
   750 => x"46415431",
   751 => x"36202020",
   752 => x"00000000",
   753 => x"46415433",
   754 => x"32202020",
   755 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;


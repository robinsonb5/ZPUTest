-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity sdbootstrap_rom is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end sdbootstrap_rom;

architecture arch of sdbootstrap_rom is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08080f4",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"97cc7383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02ec050d",
    30 => x"88bd0bff",
    31 => x"880c800b",
    32 => x"870a0cf8",
    33 => x"0883fff0",
    34 => x"900cfc08",
    35 => x"83fff094",
    36 => x"0c84eacd",
    37 => x"a8800b83",
    38 => x"fff0980c",
    39 => x"a0808790",
    40 => x"2d83ffe0",
    41 => x"8008902b",
    42 => x"70902c51",
    43 => x"5372802e",
    44 => x"81d138a0",
    45 => x"808a982d",
    46 => x"83ffe090",
    47 => x"5283fff0",
    48 => x"9051a080",
    49 => x"95a92d83",
    50 => x"ffe08008",
    51 => x"802e81b3",
    52 => x"3883ffe0",
    53 => x"90548055",
    54 => x"73708105",
    55 => x"55a08080",
    56 => x"b42d5372",
    57 => x"a02e80de",
    58 => x"3872a32e",
    59 => x"80fd3872",
    60 => x"80c72e09",
    61 => x"81068b38",
    62 => x"a0808088",
    63 => x"2da08082",
    64 => x"a204728a",
    65 => x"2e098106",
    66 => x"8b38a080",
    67 => x"80902da0",
    68 => x"8082a204",
    69 => x"7280cc2e",
    70 => x"09810686",
    71 => x"3883ffe0",
    72 => x"90547281",
    73 => x"df06f005",
    74 => x"7081ff06",
    75 => x"5153b873",
    76 => x"278938ef",
    77 => x"137081ff",
    78 => x"06515374",
    79 => x"842b7307",
    80 => x"55a08081",
    81 => x"d80472a3",
    82 => x"2ea13873",
    83 => x"70810555",
    84 => x"a08080b4",
    85 => x"2d5372a0",
    86 => x"2ef138ff",
    87 => x"14755370",
    88 => x"5254a080",
    89 => x"95a92d74",
    90 => x"870a0c73",
    91 => x"70810555",
    92 => x"a08080b4",
    93 => x"2d53728a",
    94 => x"2e098106",
    95 => x"ee38a080",
    96 => x"81d60480",
    97 => x"0b83ffe0",
    98 => x"800c0294",
    99 => x"050d0402",
   100 => x"f4050d74",
   101 => x"767181ff",
   102 => x"06c80c53",
   103 => x"5383fff0",
   104 => x"9c088538",
   105 => x"71892b52",
   106 => x"71982ac8",
   107 => x"0c71902a",
   108 => x"7081ff06",
   109 => x"c80c5171",
   110 => x"882a7081",
   111 => x"ff06c80c",
   112 => x"517181ff",
   113 => x"06c80c72",
   114 => x"902a7081",
   115 => x"ff06c80c",
   116 => x"51c80870",
   117 => x"81ff0651",
   118 => x"5182b8bf",
   119 => x"527081ff",
   120 => x"2e098106",
   121 => x"943881ff",
   122 => x"0bc80cc8",
   123 => x"087081ff",
   124 => x"06ff1454",
   125 => x"515171e5",
   126 => x"387083ff",
   127 => x"e0800c02",
   128 => x"8c050d04",
   129 => x"02fc050d",
   130 => x"81c75181",
   131 => x"ff0bc80c",
   132 => x"ff115170",
   133 => x"8025f438",
   134 => x"0284050d",
   135 => x"0402ec05",
   136 => x"0da08084",
   137 => x"842d819c",
   138 => x"9f558052",
   139 => x"87fc80f7",
   140 => x"51a08083",
   141 => x"8f2d83ff",
   142 => x"e0800890",
   143 => x"2b70902c",
   144 => x"70565153",
   145 => x"72812e09",
   146 => x"8106b338",
   147 => x"81ff0bc8",
   148 => x"0c820a52",
   149 => x"849c80e9",
   150 => x"51a08083",
   151 => x"8f2d83ff",
   152 => x"e0800890",
   153 => x"2b70902c",
   154 => x"5153728d",
   155 => x"3881ff0b",
   156 => x"c80c7353",
   157 => x"a0808587",
   158 => x"04a08084",
   159 => x"842dff15",
   160 => x"5574ffa6",
   161 => x"38745372",
   162 => x"83ffe080",
   163 => x"0c029405",
   164 => x"0d0402f0",
   165 => x"050d81ff",
   166 => x"0bc80c93",
   167 => x"54805287",
   168 => x"fc80c151",
   169 => x"a080838f",
   170 => x"2d83ffe0",
   171 => x"8008902b",
   172 => x"70902c51",
   173 => x"53728d38",
   174 => x"81ff0bc8",
   175 => x"0c8153a0",
   176 => x"8085d104",
   177 => x"a0808484",
   178 => x"2dff1454",
   179 => x"73cf3873",
   180 => x"537283ff",
   181 => x"e0800c02",
   182 => x"90050d04",
   183 => x"02f0050d",
   184 => x"a0808484",
   185 => x"2d83aa52",
   186 => x"849c80c8",
   187 => x"51a08083",
   188 => x"8f2d83ff",
   189 => x"e0800881",
   190 => x"2e098106",
   191 => x"9038cc08",
   192 => x"7083ffff",
   193 => x"06515372",
   194 => x"83aa2e99",
   195 => x"38a08085",
   196 => x"922da080",
   197 => x"869e0481",
   198 => x"54a08087",
   199 => x"85048054",
   200 => x"a0808785",
   201 => x"0481ff0b",
   202 => x"c80cb154",
   203 => x"a080849d",
   204 => x"2d83ffe0",
   205 => x"8008902b",
   206 => x"70902c51",
   207 => x"5372802e",
   208 => x"b7388052",
   209 => x"87fc80fa",
   210 => x"51a08083",
   211 => x"8f2d83ff",
   212 => x"e08008a4",
   213 => x"3881ff0b",
   214 => x"c80cc808",
   215 => x"cc087186",
   216 => x"2a708106",
   217 => x"83ffe080",
   218 => x"08535152",
   219 => x"55537280",
   220 => x"2e9338a0",
   221 => x"80869704",
   222 => x"73822eff",
   223 => x"a138ff14",
   224 => x"5473ffa8",
   225 => x"387383ff",
   226 => x"e0800c02",
   227 => x"90050d04",
   228 => x"02f4050d",
   229 => x"810b83ff",
   230 => x"f09c0cc4",
   231 => x"08708f2a",
   232 => x"70810651",
   233 => x"515372f3",
   234 => x"3872c40c",
   235 => x"a0808484",
   236 => x"2dc40870",
   237 => x"8f2a7081",
   238 => x"06515153",
   239 => x"72f33881",
   240 => x"0bc40c87",
   241 => x"53805284",
   242 => x"d480c051",
   243 => x"a080838f",
   244 => x"2d83ffe0",
   245 => x"8008812e",
   246 => x"96387282",
   247 => x"2e098106",
   248 => x"88388053",
   249 => x"a08088ad",
   250 => x"04ff1353",
   251 => x"72d738a0",
   252 => x"8085dc2d",
   253 => x"83ffe080",
   254 => x"08902b70",
   255 => x"902c83ff",
   256 => x"f09c0c53",
   257 => x"815287fc",
   258 => x"80d051a0",
   259 => x"80838f2d",
   260 => x"81ff0bc8",
   261 => x"0cc40870",
   262 => x"8f2a7081",
   263 => x"06515153",
   264 => x"72f33872",
   265 => x"c40c81ff",
   266 => x"0bc80c81",
   267 => x"537283ff",
   268 => x"e0800c02",
   269 => x"8c050d04",
   270 => x"800b83ff",
   271 => x"e0800c04",
   272 => x"02e8050d",
   273 => x"78558056",
   274 => x"c408708f",
   275 => x"2a708106",
   276 => x"51515372",
   277 => x"f3388281",
   278 => x"0bc40c81",
   279 => x"ff0bc80c",
   280 => x"775287fc",
   281 => x"80d151a0",
   282 => x"80838f2d",
   283 => x"83ffe080",
   284 => x"0880d238",
   285 => x"80dbc6df",
   286 => x"5481ff0b",
   287 => x"c80cc808",
   288 => x"7081ff06",
   289 => x"51537281",
   290 => x"fe2e0981",
   291 => x"069b3880",
   292 => x"ff54cc08",
   293 => x"75708405",
   294 => x"570cff14",
   295 => x"54738025",
   296 => x"f1388156",
   297 => x"a08089af",
   298 => x"04ff1454",
   299 => x"73cb3881",
   300 => x"ff0bc80c",
   301 => x"c408708f",
   302 => x"2a708106",
   303 => x"51515372",
   304 => x"f33872c4",
   305 => x"0c7583ff",
   306 => x"e0800c02",
   307 => x"98050d04",
   308 => x"02e8050d",
   309 => x"77797b58",
   310 => x"55558053",
   311 => x"727625ab",
   312 => x"38747081",
   313 => x"0556a080",
   314 => x"80b42d74",
   315 => x"70810556",
   316 => x"a08080b4",
   317 => x"2d525271",
   318 => x"712e8838",
   319 => x"8151a080",
   320 => x"8a8d0481",
   321 => x"1353a080",
   322 => x"89dc0480",
   323 => x"517083ff",
   324 => x"e0800c02",
   325 => x"98050d04",
   326 => x"02d8050d",
   327 => x"ff0b83ff",
   328 => x"f4c80c80",
   329 => x"0b83fff4",
   330 => x"dc0c83ff",
   331 => x"f0b45280",
   332 => x"51a08088",
   333 => x"c02d83ff",
   334 => x"e0800890",
   335 => x"2b70902c",
   336 => x"70575154",
   337 => x"73802e86",
   338 => x"d7388056",
   339 => x"810b83ff",
   340 => x"f0a80c88",
   341 => x"53a08097",
   342 => x"dc5283ff",
   343 => x"f0ea51a0",
   344 => x"8089d02d",
   345 => x"83ffe080",
   346 => x"08762e09",
   347 => x"81068b38",
   348 => x"83ffe080",
   349 => x"0883fff0",
   350 => x"a80c8853",
   351 => x"a08097e8",
   352 => x"5283fff1",
   353 => x"8651a080",
   354 => x"89d02d83",
   355 => x"ffe08008",
   356 => x"8b3883ff",
   357 => x"e0800883",
   358 => x"fff0a80c",
   359 => x"83fff0a8",
   360 => x"08802e81",
   361 => x"a03883ff",
   362 => x"f3fa0ba0",
   363 => x"8080b42d",
   364 => x"83fff3fb",
   365 => x"0ba08080",
   366 => x"b42d7198",
   367 => x"2b71902b",
   368 => x"0783fff3",
   369 => x"fc0ba080",
   370 => x"80b42d70",
   371 => x"882b7207",
   372 => x"83fff3fd",
   373 => x"0ba08080",
   374 => x"b42d7107",
   375 => x"83fff4b2",
   376 => x"0ba08080",
   377 => x"b42d83ff",
   378 => x"f4b30ba0",
   379 => x"8080b42d",
   380 => x"71882b07",
   381 => x"535f5452",
   382 => x"5a565755",
   383 => x"7381abaa",
   384 => x"2e098106",
   385 => x"93387551",
   386 => x"a08096df",
   387 => x"2d83ffe0",
   388 => x"800856a0",
   389 => x"808ca504",
   390 => x"80557382",
   391 => x"d4d52e09",
   392 => x"810684fc",
   393 => x"3883fff0",
   394 => x"b4527551",
   395 => x"a08088c0",
   396 => x"2d83ffe0",
   397 => x"8008902b",
   398 => x"70902c70",
   399 => x"57515473",
   400 => x"802e84dc",
   401 => x"388853a0",
   402 => x"8097e852",
   403 => x"83fff186",
   404 => x"51a08089",
   405 => x"d02d83ff",
   406 => x"e080088d",
   407 => x"38810b83",
   408 => x"fff4dc0c",
   409 => x"a0808d89",
   410 => x"048853a0",
   411 => x"8097dc52",
   412 => x"83fff0ea",
   413 => x"51a08089",
   414 => x"d02d8055",
   415 => x"83ffe080",
   416 => x"08752e09",
   417 => x"81068498",
   418 => x"3883fff4",
   419 => x"b20ba080",
   420 => x"80b42d54",
   421 => x"7380d52e",
   422 => x"09810680",
   423 => x"db3883ff",
   424 => x"f4b30ba0",
   425 => x"8080b42d",
   426 => x"547381aa",
   427 => x"2e098106",
   428 => x"80c63880",
   429 => x"0b83fff0",
   430 => x"b40ba080",
   431 => x"80b42d56",
   432 => x"547481e9",
   433 => x"2e833881",
   434 => x"547481eb",
   435 => x"2e8c3880",
   436 => x"5573752e",
   437 => x"09810683",
   438 => x"c73883ff",
   439 => x"f0bf0ba0",
   440 => x"8080b42d",
   441 => x"55749138",
   442 => x"83fff0c0",
   443 => x"0ba08080",
   444 => x"b42d5473",
   445 => x"822e8838",
   446 => x"8055a080",
   447 => x"91a00483",
   448 => x"fff0c10b",
   449 => x"a08080b4",
   450 => x"2d7083ff",
   451 => x"f4e40cff",
   452 => x"0583fff4",
   453 => x"d80c83ff",
   454 => x"f0c20ba0",
   455 => x"8080b42d",
   456 => x"83fff0c3",
   457 => x"0ba08080",
   458 => x"b42d5876",
   459 => x"05778280",
   460 => x"29057083",
   461 => x"fff4cc0c",
   462 => x"83fff0c4",
   463 => x"0ba08080",
   464 => x"b42d7083",
   465 => x"fff4c40c",
   466 => x"83fff4dc",
   467 => x"08595758",
   468 => x"76802e81",
   469 => x"df388853",
   470 => x"a08097e8",
   471 => x"5283fff1",
   472 => x"8651a080",
   473 => x"89d02d83",
   474 => x"ffe08008",
   475 => x"82b23883",
   476 => x"fff4e408",
   477 => x"70842b83",
   478 => x"fff4b40c",
   479 => x"7083fff4",
   480 => x"e00c83ff",
   481 => x"f0d90ba0",
   482 => x"8080b42d",
   483 => x"83fff0d8",
   484 => x"0ba08080",
   485 => x"b42d7182",
   486 => x"80290583",
   487 => x"fff0da0b",
   488 => x"a08080b4",
   489 => x"2d708480",
   490 => x"80291283",
   491 => x"fff0db0b",
   492 => x"a08080b4",
   493 => x"2d708180",
   494 => x"0a291270",
   495 => x"83fff0ac",
   496 => x"0c83fff4",
   497 => x"c4087129",
   498 => x"83fff4cc",
   499 => x"08057083",
   500 => x"fff4ec0c",
   501 => x"83fff0e1",
   502 => x"0ba08080",
   503 => x"b42d83ff",
   504 => x"f0e00ba0",
   505 => x"8080b42d",
   506 => x"71828029",
   507 => x"0583fff0",
   508 => x"e20ba080",
   509 => x"80b42d70",
   510 => x"84808029",
   511 => x"1283fff0",
   512 => x"e30ba080",
   513 => x"80b42d70",
   514 => x"982b81f0",
   515 => x"0a067205",
   516 => x"7083fff0",
   517 => x"b00cfe11",
   518 => x"7e297705",
   519 => x"83fff4d4",
   520 => x"0c525952",
   521 => x"43545e51",
   522 => x"5259525d",
   523 => x"575957a0",
   524 => x"80919e04",
   525 => x"83fff0c6",
   526 => x"0ba08080",
   527 => x"b42d83ff",
   528 => x"f0c50ba0",
   529 => x"8080b42d",
   530 => x"71828029",
   531 => x"057083ff",
   532 => x"f4b40c70",
   533 => x"a02983ff",
   534 => x"0570892a",
   535 => x"7083fff4",
   536 => x"e00c83ff",
   537 => x"f0cb0ba0",
   538 => x"8080b42d",
   539 => x"83fff0ca",
   540 => x"0ba08080",
   541 => x"b42d7182",
   542 => x"80290570",
   543 => x"83fff0ac",
   544 => x"0c7b7129",
   545 => x"1e7083ff",
   546 => x"f4d40c7d",
   547 => x"83fff0b0",
   548 => x"0c730583",
   549 => x"fff4ec0c",
   550 => x"555e5151",
   551 => x"55558155",
   552 => x"7483ffe0",
   553 => x"800c02a8",
   554 => x"050d0402",
   555 => x"e8050d77",
   556 => x"70872c71",
   557 => x"80ff0656",
   558 => x"565383ff",
   559 => x"f4dc088a",
   560 => x"3872882c",
   561 => x"7381ff06",
   562 => x"55557483",
   563 => x"fff4c808",
   564 => x"2eac3883",
   565 => x"fff0b452",
   566 => x"83fff4cc",
   567 => x"081551a0",
   568 => x"8088c02d",
   569 => x"83ffe080",
   570 => x"08902b70",
   571 => x"902c7058",
   572 => x"51537280",
   573 => x"2e80cb38",
   574 => x"7483fff4",
   575 => x"c80c83ff",
   576 => x"f4dc0880",
   577 => x"2ea03873",
   578 => x"842983ff",
   579 => x"f0b40570",
   580 => x"085253a0",
   581 => x"8096df2d",
   582 => x"83ffe080",
   583 => x"08f00a06",
   584 => x"54a08092",
   585 => x"c0047310",
   586 => x"83fff0b4",
   587 => x"0570a080",
   588 => x"809f2d52",
   589 => x"53a08097",
   590 => x"912d83ff",
   591 => x"e0800854",
   592 => x"73567583",
   593 => x"ffe0800c",
   594 => x"0298050d",
   595 => x"0402cc05",
   596 => x"0d7e605e",
   597 => x"5b8056ff",
   598 => x"0b83fff4",
   599 => x"c80c83ff",
   600 => x"f0b00883",
   601 => x"fff4d408",
   602 => x"565a83ff",
   603 => x"f4dc0876",
   604 => x"2e8e3883",
   605 => x"fff4e408",
   606 => x"842b58a0",
   607 => x"80938804",
   608 => x"83fff4e0",
   609 => x"08842b58",
   610 => x"80597878",
   611 => x"2781c938",
   612 => x"788f06a0",
   613 => x"17575473",
   614 => x"953883ff",
   615 => x"f0b45274",
   616 => x"51811555",
   617 => x"a08088c0",
   618 => x"2d83fff0",
   619 => x"b4568076",
   620 => x"a08080b4",
   621 => x"2d555773",
   622 => x"772e8338",
   623 => x"81577381",
   624 => x"e52e818c",
   625 => x"38817078",
   626 => x"06555c73",
   627 => x"802e8180",
   628 => x"388b16a0",
   629 => x"8080b42d",
   630 => x"98065776",
   631 => x"80f2388b",
   632 => x"537c5275",
   633 => x"51a08089",
   634 => x"d02d83ff",
   635 => x"e0800880",
   636 => x"df389c16",
   637 => x"0851a080",
   638 => x"96df2d83",
   639 => x"ffe08008",
   640 => x"841c0c9a",
   641 => x"16a08080",
   642 => x"9f2d51a0",
   643 => x"8097912d",
   644 => x"83ffe080",
   645 => x"0883ffe0",
   646 => x"80085555",
   647 => x"83fff4dc",
   648 => x"08802e9e",
   649 => x"389416a0",
   650 => x"80809f2d",
   651 => x"51a08097",
   652 => x"912d83ff",
   653 => x"e0800890",
   654 => x"2b83fff0",
   655 => x"0a067016",
   656 => x"51547388",
   657 => x"1c0c767b",
   658 => x"0c7b54a0",
   659 => x"80959e04",
   660 => x"811959a0",
   661 => x"80938a04",
   662 => x"83fff4dc",
   663 => x"08802ebc",
   664 => x"387951a0",
   665 => x"8091ab2d",
   666 => x"83ffe080",
   667 => x"0883ffe0",
   668 => x"800880ff",
   669 => x"fffff806",
   670 => x"555a7380",
   671 => x"fffffff8",
   672 => x"2e9a3883",
   673 => x"ffe08008",
   674 => x"fe0583ff",
   675 => x"f4e40829",
   676 => x"83fff4ec",
   677 => x"080555a0",
   678 => x"80938804",
   679 => x"80547383",
   680 => x"ffe0800c",
   681 => x"02b4050d",
   682 => x"0402e405",
   683 => x"0d797953",
   684 => x"83fff4b8",
   685 => x"5255a080",
   686 => x"92cd2d83",
   687 => x"ffe08008",
   688 => x"81ff0670",
   689 => x"55537280",
   690 => x"2e818938",
   691 => x"83fff4bc",
   692 => x"0883ff05",
   693 => x"892a5780",
   694 => x"70555675",
   695 => x"772580f2",
   696 => x"3883fff4",
   697 => x"c008fe05",
   698 => x"83fff4e4",
   699 => x"082983ff",
   700 => x"f4ec0811",
   701 => x"7583fff4",
   702 => x"d8080605",
   703 => x"76545253",
   704 => x"a08088c0",
   705 => x"2d83ffe0",
   706 => x"8008902b",
   707 => x"70902c51",
   708 => x"5372802e",
   709 => x"b6388114",
   710 => x"7083fff4",
   711 => x"d8080654",
   712 => x"54729638",
   713 => x"83fff4c0",
   714 => x"0851a080",
   715 => x"91ab2d83",
   716 => x"ffe08008",
   717 => x"83fff4c0",
   718 => x"0c848015",
   719 => x"81175755",
   720 => x"767624ff",
   721 => x"9c38a080",
   722 => x"96d20472",
   723 => x"54a08096",
   724 => x"d4048154",
   725 => x"7383ffe0",
   726 => x"800c029c",
   727 => x"050d0402",
   728 => x"f4050d74",
   729 => x"70882a83",
   730 => x"fe800670",
   731 => x"72982a07",
   732 => x"72882b87",
   733 => x"fc808006",
   734 => x"73982b81",
   735 => x"f00a0671",
   736 => x"73070783",
   737 => x"ffe0800c",
   738 => x"56515351",
   739 => x"028c050d",
   740 => x"0402f405",
   741 => x"0d029205",
   742 => x"a080809f",
   743 => x"2d70882a",
   744 => x"71882b07",
   745 => x"7083ffff",
   746 => x"0683ffe0",
   747 => x"800c5252",
   748 => x"028c050d",
   749 => x"0402f805",
   750 => x"0d737090",
   751 => x"2b71902a",
   752 => x"0783ffe0",
   753 => x"800c5202",
   754 => x"88050d04",
   755 => x"00ffffff",
   756 => x"ff00ffff",
   757 => x"ffff00ff",
   758 => x"ffffff00",
   759 => x"46415431",
   760 => x"36202020",
   761 => x"00000000",
   762 => x"46415433",
   763 => x"32202020",
   764 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;


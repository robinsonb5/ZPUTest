library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.ALL;

-- VGA controller
-- a module to handle VGA output

-- Modified for ZPU use, data bus is now 32-bits wide.

-- Self-contained, must generate timings
-- Programmable, must provide hardware registers that will respond to
-- writes.  Registers will include:  (Decode a 4k chunk)

-- 0 / 2   Framebuffer Address - hi and low
--     4   Even row modulo
--     6   Odd row modulo (allows scandoubling)

--     8  HTotal
--     A  HSize (typically 640)
--     C  HBStart
--     E  HBStop

--    10  VTotal
--    12  VSize (typically 480)
--    14  VBStart
--    16  VBStop

--    18  Control:
--     0  Visible
--     1  Resolution - high, low  - alternatively could make pixel clock programmable...
--     7  Character overlay on/off

--   Character buffer (2048 bytes)


-- Present the following signals to the SOC:
--	clk : in std_logic;
--	reset : in std_logic;

--	reg_addr_in : in std_logic_vector(10 downto 0);
--	reg_rw : std_logic;
--	reg_uds : std_logic;	-- only affects char buffer
--	reg_lds : std_logic;

	--		reqin : in std_logic;  -- now generated by VGA module
	--		data_out : out std_logic_vector(15 downto 0); -- now used internally

--		newframe : in std_logic; -- 
--		addrout : buffer std_logic_vector(23 downto 0); -- to SDRAM
--		data_in : in std_logic_vector(15 downto 0);	-- from SDRAM
--		fill : in std_logic; -- High when data is being written from SDRAM controller
--		req : buffer std_logic -- Request service from SDRAM controller

--		hsync : std_logic -- to monitor
--		vsync : std_logic -- to monitor
--		red : std_logic_vector(4 downto 0);		-- 16-bit 5-6-5 output
--		green : std_logic_vector(5 downto 0);
--		blue : std_logic_vector(4 downto 0);


-- FIXME - make address bus 32 bits wide.

entity vga_controller is
  generic(
		enable_sprite : boolean := true
	);
  port (
		clk : in std_logic;
		reset : in std_logic;

		reg_addr_in : in std_logic_vector(11 downto 0); -- from host CPU
		reg_data_in: in std_logic_vector(31 downto 0);
		reg_data_out: out std_logic_vector(15 downto 0);
		reg_rw : in std_logic;
		reg_uds : in std_logic;
		reg_lds : in std_logic;
		reg_dtack : out std_logic;	-- Needed for char ram access.
		reg_req : in std_logic;

		sdr_addrout : buffer std_logic_vector(31 downto 0); -- to SDRAM
		sdr_datain : in std_logic_vector(15 downto 0);	-- from SDRAM
		sdr_fill : in std_logic; -- High when data is being written from SDRAM controller
		sdr_req : buffer std_logic; -- Request service from SDRAM controller
		sdr_reservebank : buffer std_logic; -- Indicate to SDR controller when requests are not critical timewise
		sdr_reserveaddr : buffer std_logic_vector(31 downto 0); -- Indicate to SDR controller when requests are not critical timewise
		sdr_refresh : out std_logic;
		sdr_ack : in std_logic;

		vblank_int : out std_logic;
		hsync : out std_logic; -- to monitor
		vsync : buffer std_logic; -- to monitor
		red : out unsigned(7 downto 0);		-- Allow for 8bpp even if we
		green : out unsigned(7 downto 0);	-- only currently support 16-bit
		blue : out unsigned(7 downto 0);		-- 5-6-5 output
		vga_window : out std_logic	-- '1' during the display window
	);
end entity;
	
architecture rtl of vga_controller is
	signal vga_pointer : std_logic_vector(31 downto 0);

	signal dma_addr : std_logic_vector(31 downto 0);
	signal setaddr_vga : std_logic;
	signal setaddr_spr0 : std_logic;
	signal dma_len : unsigned(11 downto 0);
	signal setlen_vga : std_logic;
	signal setlen_spr0 : std_logic;
	signal req_vga : std_logic;
	signal req_spr0 : std_logic;
	signal data_from_dma : std_logic_vector(15 downto 0);
	signal valid_vga : std_logic;
	signal valid_spr0 : std_logic;
	
	signal framebuffer_pointer : std_logic_vector(31 downto 0) := X"00100000";
	signal hsize : unsigned(11 downto 0) := TO_UNSIGNED(640,12);
	signal htotal : unsigned(11 downto 0) := TO_UNSIGNED(800,12);
	signal hbstart : unsigned(11 downto 0) := TO_UNSIGNED(656,12);
	signal hbstop : unsigned(11 downto 0) := TO_UNSIGNED(752,12);
	signal vsize : unsigned(11 downto 0) := TO_UNSIGNED(480,12);
	signal vtotal : unsigned(11 downto 0) := TO_UNSIGNED(525,12);
	signal vbstart : unsigned(11 downto 0) := TO_UNSIGNED(500,12);
	signal vbstop : unsigned(11 downto 0) := TO_UNSIGNED(502,12);

	signal sprite0_pointer : std_logic_vector(31 downto 0) := X"00000000";
	signal sprite0_xpos : unsigned(11 downto 0);
	signal sprite0_ypos : unsigned(11 downto 0);
	signal sprite0_data : std_logic_vector(15 downto 0);
	signal sprite0_counter : unsigned(1 downto 0);

	signal sprite_col : std_logic_vector(3 downto 0);
	
	signal currentX : unsigned(11 downto 0);
	signal currentY : unsigned(11 downto 0);
	signal end_of_pixel : std_logic;
	signal vga_newframe : std_logic;
	signal vgadata : std_logic_vector(15 downto 0);

begin

	myVgaMaster : entity work.video_vga_master
		generic map (
			clkDivBits => 4
		)
		port map (
			clk => clk,
--			clkDiv => X"3",	-- 100 Mhz / (3+1) = 25 Mhz
			clkDiv => X"4",	-- 125 Mhz / (4+1) = 25 Mhz

			hSync => hsync,
			vSync => vsync,

			endOfPixel => end_of_pixel,
			endOfLine => open,
			endOfFrame => open,
			currentX => currentX,
			currentY => currentY,

			-- Setup 640x480@60hz needs ~25 Mhz
			hSyncPol => '0',
			vSyncPol => '0',
			xSize => htotal,
			ySize => vtotal,
			xSyncFr => hbstart,
			xSyncTo => hbstop,
			ySyncFr => vbstart, -- Sync pulse 2
			ySyncTo => vbstop
		);		

	mydmacache : entity work.DMACache
		port map(
			clk => clk,
			reset_n => reset,

			-- DMA addressing
			addr_in => dma_addr,
			setaddr_vga => setaddr_vga,
			setaddr_sprite0 => setaddr_spr0,
			setaddr_audio0 => '0',
			setaddr_audio1 => '0',

			-- DMA request lengths
			req_length => dma_len,
			setreqlen_vga => setlen_vga,
			setreqlen_sprite0 => setlen_spr0,
			setreqlen_audio0 => '0',
			setreqlen_audio1 => '0',

			-- Read requests
			req_vga => req_vga,
			req_sprite0 => req_spr0,
			req_audio0 => '0',
			req_audio1 => '0',

			-- DMA channel output and valid flags.
			data_out => data_from_dma,
			valid_vga => valid_vga,
			valid_sprite0 => valid_spr0,
			valid_audio0 => open,
			valid_audio1 => open,
			
			-- SDRAM interface
			sdram_addr=> sdr_addrout,
			sdram_reserveaddr(31 downto 0) => sdr_reserveaddr,
			sdram_reserve => sdr_reservebank,
			sdram_req => sdr_req,
			sdram_ack => sdr_ack,
			sdram_fill => sdr_fill,
			sdram_data => sdr_datain
		);

	-- Handle CPU access to hardware registers
	
	process(clk,reset)
	begin
		if reset='0' then
			htotal <= TO_UNSIGNED(800,12);
			vtotal <= TO_UNSIGNED(525,12);
			hbstart <= TO_UNSIGNED(656,12);
			hbstop <= TO_UNSIGNED(752,12);
			vbstart <= TO_UNSIGNED(500,12);
			vbstop <= TO_UNSIGNED(502,12);
			reg_data_out<=X"0000";
			sprite0_xpos<=X"000";
			sprite0_ypos<=X"000";
		elsif rising_edge(clk) then
			reg_dtack<='1';
			if reg_req='1' then
				case reg_addr_in is
					when X"000" =>
	--					reg_data_out<=X"00"&framebuffer_pointer(23 downto 16);
						if reg_rw='0' then
							framebuffer_pointer(31 downto 0) <= reg_data_in;
						end if;
					when X"100" =>
	--					reg_data_out<=X"00"&sprite0_pointer(23 downto 16);
						if reg_rw='0' and enable_sprite then
							sprite0_pointer(31 downto 0) <= reg_data_in;
						end if;
					when X"104" =>
						if reg_rw='0' and enable_sprite then
							sprite0_xpos <= unsigned(reg_data_in(11 downto 0));
						end if;
					when X"108" =>
						if reg_rw='0' and enable_sprite then
							sprite0_ypos <= unsigned(reg_data_in(11 downto 0));
						end if;
					when others =>
						reg_data_out<=X"0000";
				end case;
				reg_dtack<='0';
			end if;
-- FBPTH equ $0000	; Framebuffer pointer - must be 64-bit aligned.
-- FBPTL equ $0002

--     4   Even row modulo
--     6   Odd row modulo (allows scandoubling)

--     8  HTotal
--     A  HSize (typically 640)
--     C  HBStart
--     E  HBStop

--    10  VTotal
--    12  VSize (typically 480)
--    14  VBStart
--    16  VBStop

--    18  Control:
--     0  Visible
--     1  Resolution - high, low  - alternatively could make pixel clock programmable...
--     7  Character overlay on/off

-- SP0PTH equ $0100 ; Pointer to sprite 0's data - must be 64-bit aligned.
-- SP0PTL equ $0102
-- SP0XPOS	equ $0104
-- SP0YPOS equ $0106


		end if;
	end process;

	
	-- Sprite positions
	process(clk, reset, currentX, currentY)
	begin
		if rising_edge(clk) then
			req_spr0<='0';
			if enable_sprite and currentX>=sprite0_xpos and currentX-sprite0_xpos<16
						and currentY>=sprite0_ypos and currentY-sprite0_ypos<16 then	
				if end_of_pixel='1' then
					case sprite0_counter is
						when "11" =>
							sprite_col<=sprite0_data(15 downto 12);
							sprite0_counter<="10";
						when "10" =>
							sprite_col<=sprite0_data(11 downto 8);
							sprite0_counter<="01";
						when "01" =>
							sprite_col<=sprite0_data(7 downto 4);
							sprite0_counter<="00";
						when "00" =>
							sprite_col<=sprite0_data(3 downto 0);
							req_spr0<='1';
							sprite0_counter<="11";
					end case;
				end if;
			else
				sprite_col<="0000";
--				sprite0_counter<="11";
			end if;

--			Prefetch first word.
			if enable_sprite and setaddr_spr0='1' then
				req_spr0<='1';
				sprite0_counter<="11";
			end if;
			
			if enable_sprite and valid_spr0='1' then
				sprite0_data<=data_from_dma;
			end if;

		end if;
	end process;
	
	
	process(clk, reset,currentX, currentY)
	begin
		if rising_edge(clk) then
			sdr_refresh <='0';
			if end_of_pixel='1' and currentX=hsize then
				sdr_refresh<='1';
			end if;
		end if;
		
		if rising_edge(clk) then
			vblank_int<='0';
			req_vga<='0';
			vga_newframe<='0';
			setaddr_vga<='0';
			setaddr_spr0<='0';
			setlen_vga<='0';
			setlen_spr0<='0';	

			if(valid_vga='1') then
				vgadata<=data_from_dma;
			end if;

			if end_of_pixel='1' then
--				sdr_reservebank<='1';

				if currentX<640 and currentY<480 then
					vga_window<='1';
					-- Request next pixel from VGA cache
					req_vga<='1';

					if sprite_col(3)='1' then
						red <= (others => sprite_col(2));
					else
						red <= unsigned(vgadata(15 downto 11)&"000");
					end if;

					if sprite_col(3)='1' then
						green <= (others=>sprite_col(1));
					else
						green <= unsigned(vgadata(10 downto 5)&"00");
					end if;

					if sprite_col(3)='1' then
						blue <= (others=>sprite_col(0));
					else
						blue <= unsigned(vgadata(4 downto 0)&"000");
					end if;

				else
					vga_window<='0';
					
					-- New frame...
					if currentY=vsize and currentX=0 then
						vblank_int<='1';
					end if;

					-- Last line of VBLANK - update DMA pointers
					if currentY=vtotal then
							if currentX=0 then
								dma_addr<=framebuffer_pointer;
								setaddr_vga<='1';
							elsif currentX=1 then
								dma_addr<=sprite0_pointer;
								setaddr_spr0<='1';
							end if;
					end if;
					
--					if currentX>(hsize+12) and currentX<(htotal - 4) then	-- Signal to SDRAM controller that we're
					if currentX=(htotal - 20) then	-- Signal to SDRAM controller that we're
						dma_len<=TO_UNSIGNED(640,12);
						setlen_vga<='1';
--						sdr_reservebank<='0'; -- in blank areas, so there's no need to keep slot 2 off the next bank.
					elsif enable_sprite and currentX=(htotal - 19) then
						dma_len<=TO_UNSIGNED(4,12);
						setlen_spr0<='1';
					end if;
				end if;
			end if;
		end if;
	end process;
		
end architecture;
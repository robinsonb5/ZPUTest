     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80c1d00c",
     3 => x"3a0b0b0b",
     4 => x"aaa30400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"8f040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bb5",
   162 => x"a4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f7040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"df040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80c1cc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"83e13fac",
   257 => x"f43f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104b0",
   280 => x"08b408b8",
   281 => x"087575a4",
   282 => x"c92d5050",
   283 => x"b00856b8",
   284 => x"0cb40cb0",
   285 => x"0c5104b0",
   286 => x"08b408b8",
   287 => x"087575a3",
   288 => x"972d5050",
   289 => x"b00856b8",
   290 => x"0cb40cb0",
   291 => x"0c5104b0",
   292 => x"08b408b8",
   293 => x"08aaea2d",
   294 => x"b80cb40c",
   295 => x"b00c04fe",
   296 => x"3d0d0b0b",
   297 => x"80c8fc08",
   298 => x"53841308",
   299 => x"70882a70",
   300 => x"81065152",
   301 => x"5270802e",
   302 => x"f0387181",
   303 => x"ff06b00c",
   304 => x"843d0d04",
   305 => x"ff3d0d0b",
   306 => x"0b80c8fc",
   307 => x"08527108",
   308 => x"70882a81",
   309 => x"32708106",
   310 => x"51515170",
   311 => x"f1387372",
   312 => x"0c833d0d",
   313 => x"0480c1cc",
   314 => x"08802ea4",
   315 => x"3880c1d0",
   316 => x"08822ebd",
   317 => x"38838080",
   318 => x"0b0b0b80",
   319 => x"c8fc0c82",
   320 => x"a0800b80",
   321 => x"c9800c82",
   322 => x"90800b80",
   323 => x"c9840c04",
   324 => x"f8808080",
   325 => x"a40b0b0b",
   326 => x"80c8fc0c",
   327 => x"f8808082",
   328 => x"800b80c9",
   329 => x"800cf880",
   330 => x"8084800b",
   331 => x"80c9840c",
   332 => x"0480c0a8",
   333 => x"808c0b0b",
   334 => x"0b80c8fc",
   335 => x"0c80c0a8",
   336 => x"80940b80",
   337 => x"c9800cb5",
   338 => x"b40b80c9",
   339 => x"840c04f2",
   340 => x"3d0d6080",
   341 => x"c9800856",
   342 => x"5d82750c",
   343 => x"8059805a",
   344 => x"800b8f3d",
   345 => x"5d5b7a10",
   346 => x"10157008",
   347 => x"7108719f",
   348 => x"2c7e852b",
   349 => x"5855557d",
   350 => x"53595796",
   351 => x"a43f7d7f",
   352 => x"7a72077c",
   353 => x"72077171",
   354 => x"60810541",
   355 => x"5f5d5b59",
   356 => x"5755817b",
   357 => x"278f3876",
   358 => x"7d0c7784",
   359 => x"1e0c7cb0",
   360 => x"0c903d0d",
   361 => x"0480c980",
   362 => x"0855ffba",
   363 => x"39ff3d0d",
   364 => x"80c98833",
   365 => x"5170a738",
   366 => x"80c1d808",
   367 => x"70085252",
   368 => x"70802e94",
   369 => x"38841280",
   370 => x"c1d80c70",
   371 => x"2d80c1d8",
   372 => x"08700852",
   373 => x"5270ee38",
   374 => x"810b80c9",
   375 => x"8834833d",
   376 => x"0d040480",
   377 => x"3d0d0b0b",
   378 => x"80c8f808",
   379 => x"802e8e38",
   380 => x"0b0b0b0b",
   381 => x"800b802e",
   382 => x"09810685",
   383 => x"38823d0d",
   384 => x"040b0b80",
   385 => x"c8f8510b",
   386 => x"0b0bf3f4",
   387 => x"3f823d0d",
   388 => x"0404c008",
   389 => x"b00c0402",
   390 => x"fc050d80",
   391 => x"c10b8198",
   392 => x"ec34800b",
   393 => x"819b840c",
   394 => x"70b00c02",
   395 => x"84050d04",
   396 => x"02f8050d",
   397 => x"800b8198",
   398 => x"ec335252",
   399 => x"7080c12e",
   400 => x"9a387181",
   401 => x"9b840807",
   402 => x"819b840c",
   403 => x"80c20b81",
   404 => x"98f03470",
   405 => x"b00c0288",
   406 => x"050d0481",
   407 => x"0b819b84",
   408 => x"0807819b",
   409 => x"840c80c2",
   410 => x"0b8198f0",
   411 => x"3470b00c",
   412 => x"0288050d",
   413 => x"0402f005",
   414 => x"0d757008",
   415 => x"8a055353",
   416 => x"8198ec33",
   417 => x"517080c1",
   418 => x"2e8c3873",
   419 => x"f33870b0",
   420 => x"0c029005",
   421 => x"0d04ff12",
   422 => x"708198e8",
   423 => x"0831740c",
   424 => x"b00c0290",
   425 => x"050d0402",
   426 => x"ec050d81",
   427 => x"99940855",
   428 => x"74802e8c",
   429 => x"38767508",
   430 => x"710c8199",
   431 => x"94085654",
   432 => x"8c155381",
   433 => x"98e80852",
   434 => x"8a519ae1",
   435 => x"2d73b00c",
   436 => x"0294050d",
   437 => x"0402e805",
   438 => x"0d777008",
   439 => x"5656b053",
   440 => x"81999408",
   441 => x"527451a7",
   442 => x"f52d850b",
   443 => x"8c170c85",
   444 => x"0b8c160c",
   445 => x"7508750c",
   446 => x"81999408",
   447 => x"5473802e",
   448 => x"8a387308",
   449 => x"750c8199",
   450 => x"9408548c",
   451 => x"14538198",
   452 => x"e808528a",
   453 => x"519ae12d",
   454 => x"841508ae",
   455 => x"38860b8c",
   456 => x"160c8815",
   457 => x"52881608",
   458 => x"5199fb2d",
   459 => x"81999408",
   460 => x"7008760c",
   461 => x"548c1570",
   462 => x"54548a52",
   463 => x"7308519a",
   464 => x"e12d73b0",
   465 => x"0c029805",
   466 => x"0d047508",
   467 => x"54b05373",
   468 => x"527551a7",
   469 => x"f52d73b0",
   470 => x"0c029805",
   471 => x"0d0402c8",
   472 => x"050d88bd",
   473 => x"0bff880c",
   474 => x"8198800b",
   475 => x"8198b40c",
   476 => x"8198b80b",
   477 => x"8199940c",
   478 => x"8198800b",
   479 => x"8198b80c",
   480 => x"800b8198",
   481 => x"b80b8405",
   482 => x"0c820b81",
   483 => x"98b80b88",
   484 => x"050ca80b",
   485 => x"8198b80b",
   486 => x"8c050c9f",
   487 => x"53b5b852",
   488 => x"8198c851",
   489 => x"a7f52d9f",
   490 => x"53b5d852",
   491 => x"819ae451",
   492 => x"a7f52d8a",
   493 => x"0b80d6cc",
   494 => x"0cbffc51",
   495 => x"9e962db5",
   496 => x"f8519e96",
   497 => x"2dbffc51",
   498 => x"9e962d80",
   499 => x"c1e00880",
   500 => x"2e888d38",
   501 => x"b6a8519e",
   502 => x"962dbffc",
   503 => x"519e962d",
   504 => x"80c1dc08",
   505 => x"52b6d451",
   506 => x"9e962dc0",
   507 => x"0880c9ec",
   508 => x"0c815880",
   509 => x"0b80c1dc",
   510 => x"082582e6",
   511 => x"3802ac05",
   512 => x"5b80c10b",
   513 => x"8198ec34",
   514 => x"810b819b",
   515 => x"840c80c2",
   516 => x"0b8198f0",
   517 => x"34825c83",
   518 => x"5a9f53b7",
   519 => x"84528198",
   520 => x"f451a7f5",
   521 => x"2d815d80",
   522 => x"0b8198f4",
   523 => x"53819ae4",
   524 => x"52559cc4",
   525 => x"2db00875",
   526 => x"2e098106",
   527 => x"83388155",
   528 => x"74819b84",
   529 => x"0c7b7057",
   530 => x"55748325",
   531 => x"a2387482",
   532 => x"2b7605fd",
   533 => x"055e02b8",
   534 => x"05fc0553",
   535 => x"83527551",
   536 => x"9ae12d81",
   537 => x"1c705d70",
   538 => x"57558375",
   539 => x"24e0387d",
   540 => x"54745380",
   541 => x"c9f05281",
   542 => x"999c519a",
   543 => x"f32d8199",
   544 => x"94087008",
   545 => x"5757b053",
   546 => x"76527551",
   547 => x"a7f52d85",
   548 => x"0b8c180c",
   549 => x"850b8c17",
   550 => x"0c760876",
   551 => x"0c819994",
   552 => x"08557480",
   553 => x"2e8a3874",
   554 => x"08760c81",
   555 => x"99940855",
   556 => x"8c155381",
   557 => x"98e80852",
   558 => x"8a519ae1",
   559 => x"2d841608",
   560 => x"87f03886",
   561 => x"0b8c170c",
   562 => x"88165288",
   563 => x"17085199",
   564 => x"fb2d8199",
   565 => x"94087008",
   566 => x"770c558c",
   567 => x"16705457",
   568 => x"8a527608",
   569 => x"519ae12d",
   570 => x"80c10b81",
   571 => x"98f03356",
   572 => x"56757526",
   573 => x"a23880c3",
   574 => x"5275519c",
   575 => x"972db008",
   576 => x"7d2e86ff",
   577 => x"38811670",
   578 => x"81ff0681",
   579 => x"98f03357",
   580 => x"57577476",
   581 => x"27e0387b",
   582 => x"527951a7",
   583 => x"932db008",
   584 => x"7e7054b0",
   585 => x"0853565a",
   586 => x"a3972db0",
   587 => x"085c7975",
   588 => x"3170832b",
   589 => x"707231b0",
   590 => x"0831b008",
   591 => x"8a058198",
   592 => x"ec338198",
   593 => x"e8085b54",
   594 => x"525c5657",
   595 => x"7680c12e",
   596 => x"86f83878",
   597 => x"f7388118",
   598 => x"5880c1dc",
   599 => x"087825fd",
   600 => x"a038c008",
   601 => x"8198b00c",
   602 => x"b7a4519e",
   603 => x"962dbffc",
   604 => x"519e962d",
   605 => x"b7b4519e",
   606 => x"962dbffc",
   607 => x"519e962d",
   608 => x"8198e808",
   609 => x"52b7ec51",
   610 => x"9e962d85",
   611 => x"52b88851",
   612 => x"9e962d81",
   613 => x"9b840852",
   614 => x"b8a4519e",
   615 => x"962d8152",
   616 => x"b888519e",
   617 => x"962d8198",
   618 => x"ec3352b8",
   619 => x"c0519e96",
   620 => x"2d80c152",
   621 => x"b8dc519e",
   622 => x"962d8198",
   623 => x"f03352b8",
   624 => x"f8519e96",
   625 => x"2d80c252",
   626 => x"b8dc519e",
   627 => x"962d8199",
   628 => x"bc0852b9",
   629 => x"94519e96",
   630 => x"2d8752b8",
   631 => x"88519e96",
   632 => x"2d80d6cc",
   633 => x"0852b9b0",
   634 => x"519e962d",
   635 => x"b9cc519e",
   636 => x"962db9f8",
   637 => x"519e962d",
   638 => x"81999408",
   639 => x"70085356",
   640 => x"ba84519e",
   641 => x"962dbaa0",
   642 => x"519e962d",
   643 => x"81999408",
   644 => x"84110853",
   645 => x"5bbad451",
   646 => x"9e962d80",
   647 => x"52b88851",
   648 => x"9e962d81",
   649 => x"99940888",
   650 => x"11085358",
   651 => x"baf0519e",
   652 => x"962d8252",
   653 => x"b888519e",
   654 => x"962d8199",
   655 => x"94088c11",
   656 => x"085359bb",
   657 => x"8c519e96",
   658 => x"2d9152b8",
   659 => x"88519e96",
   660 => x"2d819994",
   661 => x"08900552",
   662 => x"bba8519e",
   663 => x"962dbbc4",
   664 => x"519e962d",
   665 => x"bbfc519e",
   666 => x"962d8198",
   667 => x"b4087008",
   668 => x"5355ba84",
   669 => x"519e962d",
   670 => x"bc90519e",
   671 => x"962d8198",
   672 => x"b4088411",
   673 => x"085357ba",
   674 => x"d4519e96",
   675 => x"2d8052b8",
   676 => x"88519e96",
   677 => x"2d8198b4",
   678 => x"08881108",
   679 => x"5356baf0",
   680 => x"519e962d",
   681 => x"8152b888",
   682 => x"519e962d",
   683 => x"8198b408",
   684 => x"8c110853",
   685 => x"5bbb8c51",
   686 => x"9e962d92",
   687 => x"52b88851",
   688 => x"9e962d81",
   689 => x"98b40890",
   690 => x"0552bba8",
   691 => x"519e962d",
   692 => x"bbc4519e",
   693 => x"962d7b52",
   694 => x"bcd0519e",
   695 => x"962d8552",
   696 => x"b888519e",
   697 => x"962d7952",
   698 => x"bcec519e",
   699 => x"962d8d52",
   700 => x"b888519e",
   701 => x"962d7d52",
   702 => x"bd88519e",
   703 => x"962d8752",
   704 => x"b888519e",
   705 => x"962d7c52",
   706 => x"bda4519e",
   707 => x"962d8152",
   708 => x"b888519e",
   709 => x"962d819a",
   710 => x"e452bdc0",
   711 => x"519e962d",
   712 => x"bddc519e",
   713 => x"962d8198",
   714 => x"f452be94",
   715 => x"519e962d",
   716 => x"beb0519e",
   717 => x"962dbffc",
   718 => x"519e962d",
   719 => x"8198b008",
   720 => x"80c9ec08",
   721 => x"317080c9",
   722 => x"e80c52be",
   723 => x"e8519e96",
   724 => x"2d80c9e8",
   725 => x"085680f7",
   726 => x"7625818b",
   727 => x"3887e852",
   728 => x"7551a793",
   729 => x"2d80c1dc",
   730 => x"087053b0",
   731 => x"08525aa3",
   732 => x"972db008",
   733 => x"80c9e00c",
   734 => x"87e85279",
   735 => x"51a7932d",
   736 => x"7552b008",
   737 => x"51a3972d",
   738 => x"b00880c9",
   739 => x"e40c84b9",
   740 => x"527951a7",
   741 => x"932d7552",
   742 => x"b00851a3",
   743 => x"972db008",
   744 => x"8199980c",
   745 => x"bef8519e",
   746 => x"962d80c9",
   747 => x"e00852bf",
   748 => x"a8519e96",
   749 => x"2dbfb051",
   750 => x"9e962d80",
   751 => x"c9e40852",
   752 => x"bfa8519e",
   753 => x"962d8199",
   754 => x"980852bf",
   755 => x"e0519e96",
   756 => x"2dbffc51",
   757 => x"9e962d80",
   758 => x"0bb00c02",
   759 => x"b8050d04",
   760 => x"80c08051",
   761 => x"8fd70480",
   762 => x"c0b0519e",
   763 => x"962d80c0",
   764 => x"e8519e96",
   765 => x"2dbffc51",
   766 => x"9e962d80",
   767 => x"c9e80856",
   768 => x"87e85275",
   769 => x"51a7932d",
   770 => x"80c1dc08",
   771 => x"7053b008",
   772 => x"525aa397",
   773 => x"2db00880",
   774 => x"c9e00c87",
   775 => x"e8527951",
   776 => x"a7932d75",
   777 => x"52b00851",
   778 => x"a3972db0",
   779 => x"0880c9e4",
   780 => x"0c84b952",
   781 => x"7951a793",
   782 => x"2d7552b0",
   783 => x"0851a397",
   784 => x"2db00881",
   785 => x"99980cbe",
   786 => x"f8519e96",
   787 => x"2d80c9e0",
   788 => x"0852bfa8",
   789 => x"519e962d",
   790 => x"bfb0519e",
   791 => x"962d80c9",
   792 => x"e40852bf",
   793 => x"a8519e96",
   794 => x"2d819998",
   795 => x"0852bfe0",
   796 => x"519e962d",
   797 => x"bffc519e",
   798 => x"962d800b",
   799 => x"b00c02b8",
   800 => x"050d0402",
   801 => x"b805f805",
   802 => x"52805199",
   803 => x"fb2d9f53",
   804 => x"80c18852",
   805 => x"8198f451",
   806 => x"a7f52d77",
   807 => x"788198e8",
   808 => x"0c811770",
   809 => x"81ff0681",
   810 => x"98f03358",
   811 => x"58585a92",
   812 => x"92047608",
   813 => x"56b05375",
   814 => x"527651a7",
   815 => x"f52d80c1",
   816 => x"0b8198f0",
   817 => x"33565691",
   818 => x"f104ff15",
   819 => x"7077317c",
   820 => x"0c59800b",
   821 => x"81195959",
   822 => x"80c1dc08",
   823 => x"7825f6a1",
   824 => x"3892e204",
   825 => x"02f8050d",
   826 => x"73823270",
   827 => x"30707207",
   828 => x"8025b00c",
   829 => x"52520288",
   830 => x"050d0402",
   831 => x"f4050d74",
   832 => x"76715354",
   833 => x"5271822e",
   834 => x"83388351",
   835 => x"71812e9b",
   836 => x"38817226",
   837 => x"a0387182",
   838 => x"2ebc3871",
   839 => x"842eac38",
   840 => x"70730c70",
   841 => x"b00c028c",
   842 => x"050d0480",
   843 => x"e40b8198",
   844 => x"e808258c",
   845 => x"3880730c",
   846 => x"70b00c02",
   847 => x"8c050d04",
   848 => x"83730c70",
   849 => x"b00c028c",
   850 => x"050d0482",
   851 => x"730c70b0",
   852 => x"0c028c05",
   853 => x"0d048173",
   854 => x"0c70b00c",
   855 => x"028c050d",
   856 => x"0402fc05",
   857 => x"0d747414",
   858 => x"8205710c",
   859 => x"b00c0284",
   860 => x"050d0402",
   861 => x"d8050d7b",
   862 => x"7d7f6185",
   863 => x"1270822b",
   864 => x"75117074",
   865 => x"71708405",
   866 => x"530c5a5a",
   867 => x"5d5b760c",
   868 => x"7980f818",
   869 => x"0c798612",
   870 => x"5257585b",
   871 => x"59757725",
   872 => x"ac3881cc",
   873 => x"527651a7",
   874 => x"932db008",
   875 => x"1afc1108",
   876 => x"8105fc12",
   877 => x"0c791970",
   878 => x"089fa013",
   879 => x"0c5b5785",
   880 => x"0b8198e8",
   881 => x"0c76b00c",
   882 => x"02a8050d",
   883 => x"04b25276",
   884 => x"51a7932d",
   885 => x"b0081782",
   886 => x"2b7a1151",
   887 => x"53767370",
   888 => x"8405550c",
   889 => x"81145475",
   890 => x"7425f238",
   891 => x"81cc5276",
   892 => x"51a7932d",
   893 => x"b0081afc",
   894 => x"11088105",
   895 => x"fc120c79",
   896 => x"1970089f",
   897 => x"a0130c5b",
   898 => x"57850b81",
   899 => x"98e80c76",
   900 => x"b00c02a8",
   901 => x"050d0402",
   902 => x"f4050d02",
   903 => x"93053351",
   904 => x"80028405",
   905 => x"97053354",
   906 => x"5270732e",
   907 => x"893871b0",
   908 => x"0c028c05",
   909 => x"0d047081",
   910 => x"98ec3481",
   911 => x"0bb00c02",
   912 => x"8c050d04",
   913 => x"02dc050d",
   914 => x"7a7c5956",
   915 => x"820b8319",
   916 => x"55557416",
   917 => x"70337533",
   918 => x"5b515372",
   919 => x"792e80c7",
   920 => x"3880c10b",
   921 => x"81168116",
   922 => x"56565782",
   923 => x"7525e338",
   924 => x"ffa91770",
   925 => x"81ff0655",
   926 => x"59738226",
   927 => x"83388755",
   928 => x"81537680",
   929 => x"d22e9838",
   930 => x"77527551",
   931 => x"a98e2d80",
   932 => x"5372b008",
   933 => x"25893887",
   934 => x"158198e8",
   935 => x"0c815372",
   936 => x"b00c02a4",
   937 => x"050d0472",
   938 => x"8198ec34",
   939 => x"827525ff",
   940 => x"a1389cf0",
   941 => x"0402f405",
   942 => x"0d747033",
   943 => x"7081ff06",
   944 => x"53535370",
   945 => x"802ea738",
   946 => x"ff840870",
   947 => x"882a7081",
   948 => x"06515151",
   949 => x"70802ef0",
   950 => x"387181ff",
   951 => x"06811454",
   952 => x"ff840c72",
   953 => x"337081ff",
   954 => x"06525270",
   955 => x"db38028c",
   956 => x"050d0402",
   957 => x"f8050d02",
   958 => x"8f053352",
   959 => x"ff840870",
   960 => x"882a7081",
   961 => x"06515151",
   962 => x"70802ef0",
   963 => x"3871ff84",
   964 => x"0c028805",
   965 => x"0d0402d0",
   966 => x"050d02b4",
   967 => x"05707084",
   968 => x"0552089d",
   969 => x"f35b555b",
   970 => x"80747081",
   971 => x"05563375",
   972 => x"5a545772",
   973 => x"772ebe38",
   974 => x"72a52e09",
   975 => x"810680c6",
   976 => x"38777081",
   977 => x"05593353",
   978 => x"7280e42e",
   979 => x"81b83872",
   980 => x"80e42480",
   981 => x"c8387280",
   982 => x"e32ea238",
   983 => x"8052a551",
   984 => x"782d8052",
   985 => x"7251782d",
   986 => x"82175777",
   987 => x"70810559",
   988 => x"335372c4",
   989 => x"3876b00c",
   990 => x"02b0050d",
   991 => x"047a841c",
   992 => x"83123355",
   993 => x"5c568052",
   994 => x"7251782d",
   995 => x"81177870",
   996 => x"81055a33",
   997 => x"545772ff",
   998 => x"9f389ef5",
   999 => x"047280f3",
  1000 => x"2e098106",
  1001 => x"ffb6387a",
  1002 => x"841c7108",
  1003 => x"585c5480",
  1004 => x"76335b55",
  1005 => x"79752e8d",
  1006 => x"38811570",
  1007 => x"17703355",
  1008 => x"5b5572f5",
  1009 => x"38ff1554",
  1010 => x"807525ff",
  1011 => x"9e387570",
  1012 => x"81055733",
  1013 => x"53805272",
  1014 => x"51782d81",
  1015 => x"1774ff16",
  1016 => x"56565780",
  1017 => x"7525ff83",
  1018 => x"38757081",
  1019 => x"05573353",
  1020 => x"80527251",
  1021 => x"782d8117",
  1022 => x"74ff1656",
  1023 => x"56577480",
  1024 => x"24cc389e",
  1025 => x"eb047a84",
  1026 => x"1c710881",
  1027 => x"9b980b80",
  1028 => x"c98c545d",
  1029 => x"565c5580",
  1030 => x"5673762e",
  1031 => x"098106b8",
  1032 => x"38b00b80",
  1033 => x"c98c3481",
  1034 => x"1553ff13",
  1035 => x"5372337a",
  1036 => x"7081055c",
  1037 => x"34811656",
  1038 => x"7280c98c",
  1039 => x"2e098106",
  1040 => x"e938807a",
  1041 => x"3475819b",
  1042 => x"980bff12",
  1043 => x"56575574",
  1044 => x"8024fefa",
  1045 => x"389eeb04",
  1046 => x"738f0680",
  1047 => x"c1a80553",
  1048 => x"72337570",
  1049 => x"81055734",
  1050 => x"73842a54",
  1051 => x"73ea3880",
  1052 => x"f8757081",
  1053 => x"05573474",
  1054 => x"53b07370",
  1055 => x"81055534",
  1056 => x"7280c98c",
  1057 => x"2effbb38",
  1058 => x"ff135372",
  1059 => x"337a7081",
  1060 => x"055c3481",
  1061 => x"16567280",
  1062 => x"c98c2eff",
  1063 => x"a538a0aa",
  1064 => x"04bc0802",
  1065 => x"bc0cf53d",
  1066 => x"0dbc0894",
  1067 => x"05089d38",
  1068 => x"bc088c05",
  1069 => x"08bc0890",
  1070 => x"0508bc08",
  1071 => x"88050858",
  1072 => x"56547376",
  1073 => x"0c748417",
  1074 => x"0c81bf39",
  1075 => x"800bbc08",
  1076 => x"f0050c80",
  1077 => x"0bbc08f4",
  1078 => x"050cbc08",
  1079 => x"8c0508bc",
  1080 => x"08900508",
  1081 => x"565473bc",
  1082 => x"08f0050c",
  1083 => x"74bc08f4",
  1084 => x"050cbc08",
  1085 => x"f805bc08",
  1086 => x"f0055656",
  1087 => x"88705475",
  1088 => x"53765254",
  1089 => x"85ef3fa0",
  1090 => x"0bbc0894",
  1091 => x"050831bc",
  1092 => x"08ec050c",
  1093 => x"bc08ec05",
  1094 => x"0880249d",
  1095 => x"38800bbc",
  1096 => x"08f4050c",
  1097 => x"bc08ec05",
  1098 => x"0830bc08",
  1099 => x"fc050871",
  1100 => x"2bbc08f0",
  1101 => x"050c54b9",
  1102 => x"39bc08fc",
  1103 => x"0508bc08",
  1104 => x"ec05082a",
  1105 => x"bc08e805",
  1106 => x"0cbc08fc",
  1107 => x"0508bc08",
  1108 => x"9405082b",
  1109 => x"bc08f405",
  1110 => x"0cbc08f8",
  1111 => x"0508bc08",
  1112 => x"9405082b",
  1113 => x"70bc08e8",
  1114 => x"050807bc",
  1115 => x"08f0050c",
  1116 => x"54bc08f0",
  1117 => x"0508bc08",
  1118 => x"f40508bc",
  1119 => x"08880508",
  1120 => x"58565473",
  1121 => x"760c7484",
  1122 => x"170cbc08",
  1123 => x"880508b0",
  1124 => x"0c8d3d0d",
  1125 => x"bc0c04bc",
  1126 => x"0802bc0c",
  1127 => x"f93d0d80",
  1128 => x"0bbc08fc",
  1129 => x"050cbc08",
  1130 => x"88050880",
  1131 => x"25ab38bc",
  1132 => x"08880508",
  1133 => x"30bc0888",
  1134 => x"050c800b",
  1135 => x"bc08f405",
  1136 => x"0cbc08fc",
  1137 => x"05088838",
  1138 => x"810bbc08",
  1139 => x"f4050cbc",
  1140 => x"08f40508",
  1141 => x"bc08fc05",
  1142 => x"0cbc088c",
  1143 => x"05088025",
  1144 => x"ab38bc08",
  1145 => x"8c050830",
  1146 => x"bc088c05",
  1147 => x"0c800bbc",
  1148 => x"08f0050c",
  1149 => x"bc08fc05",
  1150 => x"08883881",
  1151 => x"0bbc08f0",
  1152 => x"050cbc08",
  1153 => x"f00508bc",
  1154 => x"08fc050c",
  1155 => x"8053bc08",
  1156 => x"8c050852",
  1157 => x"bc088805",
  1158 => x"085181a7",
  1159 => x"3fb00870",
  1160 => x"bc08f805",
  1161 => x"0c54bc08",
  1162 => x"fc050880",
  1163 => x"2e8c38bc",
  1164 => x"08f80508",
  1165 => x"30bc08f8",
  1166 => x"050cbc08",
  1167 => x"f8050870",
  1168 => x"b00c5489",
  1169 => x"3d0dbc0c",
  1170 => x"04bc0802",
  1171 => x"bc0cfb3d",
  1172 => x"0d800bbc",
  1173 => x"08fc050c",
  1174 => x"bc088805",
  1175 => x"08802593",
  1176 => x"38bc0888",
  1177 => x"050830bc",
  1178 => x"0888050c",
  1179 => x"810bbc08",
  1180 => x"fc050cbc",
  1181 => x"088c0508",
  1182 => x"80258c38",
  1183 => x"bc088c05",
  1184 => x"0830bc08",
  1185 => x"8c050c81",
  1186 => x"53bc088c",
  1187 => x"050852bc",
  1188 => x"08880508",
  1189 => x"51ad3fb0",
  1190 => x"0870bc08",
  1191 => x"f8050c54",
  1192 => x"bc08fc05",
  1193 => x"08802e8c",
  1194 => x"38bc08f8",
  1195 => x"050830bc",
  1196 => x"08f8050c",
  1197 => x"bc08f805",
  1198 => x"0870b00c",
  1199 => x"54873d0d",
  1200 => x"bc0c04bc",
  1201 => x"0802bc0c",
  1202 => x"fd3d0d81",
  1203 => x"0bbc08fc",
  1204 => x"050c800b",
  1205 => x"bc08f805",
  1206 => x"0cbc088c",
  1207 => x"0508bc08",
  1208 => x"88050827",
  1209 => x"ac38bc08",
  1210 => x"fc050880",
  1211 => x"2ea33880",
  1212 => x"0bbc088c",
  1213 => x"05082499",
  1214 => x"38bc088c",
  1215 => x"050810bc",
  1216 => x"088c050c",
  1217 => x"bc08fc05",
  1218 => x"0810bc08",
  1219 => x"fc050cc9",
  1220 => x"39bc08fc",
  1221 => x"0508802e",
  1222 => x"80c938bc",
  1223 => x"088c0508",
  1224 => x"bc088805",
  1225 => x"0826a138",
  1226 => x"bc088805",
  1227 => x"08bc088c",
  1228 => x"050831bc",
  1229 => x"0888050c",
  1230 => x"bc08f805",
  1231 => x"08bc08fc",
  1232 => x"050807bc",
  1233 => x"08f8050c",
  1234 => x"bc08fc05",
  1235 => x"08812abc",
  1236 => x"08fc050c",
  1237 => x"bc088c05",
  1238 => x"08812abc",
  1239 => x"088c050c",
  1240 => x"ffaf39bc",
  1241 => x"08900508",
  1242 => x"802e8f38",
  1243 => x"bc088805",
  1244 => x"0870bc08",
  1245 => x"f4050c51",
  1246 => x"8d39bc08",
  1247 => x"f8050870",
  1248 => x"bc08f405",
  1249 => x"0c51bc08",
  1250 => x"f40508b0",
  1251 => x"0c853d0d",
  1252 => x"bc0c04bc",
  1253 => x"0802bc0c",
  1254 => x"ff3d0d80",
  1255 => x"0bbc08fc",
  1256 => x"050cbc08",
  1257 => x"88050881",
  1258 => x"06ff1170",
  1259 => x"0970bc08",
  1260 => x"8c050806",
  1261 => x"bc08fc05",
  1262 => x"0811bc08",
  1263 => x"fc050cbc",
  1264 => x"08880508",
  1265 => x"812abc08",
  1266 => x"88050cbc",
  1267 => x"088c0508",
  1268 => x"10bc088c",
  1269 => x"050c5151",
  1270 => x"5151bc08",
  1271 => x"88050880",
  1272 => x"2e8438ff",
  1273 => x"bd39bc08",
  1274 => x"fc050870",
  1275 => x"b00c5183",
  1276 => x"3d0dbc0c",
  1277 => x"04fc3d0d",
  1278 => x"7670797b",
  1279 => x"55555555",
  1280 => x"8f72278c",
  1281 => x"38727507",
  1282 => x"83065170",
  1283 => x"802ea738",
  1284 => x"ff125271",
  1285 => x"ff2e9838",
  1286 => x"72708105",
  1287 => x"54337470",
  1288 => x"81055634",
  1289 => x"ff125271",
  1290 => x"ff2e0981",
  1291 => x"06ea3874",
  1292 => x"b00c863d",
  1293 => x"0d047451",
  1294 => x"72708405",
  1295 => x"54087170",
  1296 => x"8405530c",
  1297 => x"72708405",
  1298 => x"54087170",
  1299 => x"8405530c",
  1300 => x"72708405",
  1301 => x"54087170",
  1302 => x"8405530c",
  1303 => x"72708405",
  1304 => x"54087170",
  1305 => x"8405530c",
  1306 => x"f0125271",
  1307 => x"8f26c938",
  1308 => x"83722795",
  1309 => x"38727084",
  1310 => x"05540871",
  1311 => x"70840553",
  1312 => x"0cfc1252",
  1313 => x"718326ed",
  1314 => x"387054ff",
  1315 => x"8339fb3d",
  1316 => x"0d777970",
  1317 => x"72078306",
  1318 => x"53545270",
  1319 => x"93387173",
  1320 => x"73085456",
  1321 => x"54717308",
  1322 => x"2e80c438",
  1323 => x"73755452",
  1324 => x"71337081",
  1325 => x"ff065254",
  1326 => x"70802e9d",
  1327 => x"38723355",
  1328 => x"70752e09",
  1329 => x"81069538",
  1330 => x"81128114",
  1331 => x"71337081",
  1332 => x"ff065456",
  1333 => x"545270e5",
  1334 => x"38723355",
  1335 => x"7381ff06",
  1336 => x"7581ff06",
  1337 => x"717131b0",
  1338 => x"0c525287",
  1339 => x"3d0d0471",
  1340 => x"0970f7fb",
  1341 => x"fdff1406",
  1342 => x"70f88482",
  1343 => x"81800651",
  1344 => x"51517097",
  1345 => x"38841484",
  1346 => x"16710854",
  1347 => x"56547175",
  1348 => x"082edc38",
  1349 => x"73755452",
  1350 => x"ff963980",
  1351 => x"0bb00c87",
  1352 => x"3d0d04fd",
  1353 => x"3d0d800b",
  1354 => x"80c1d008",
  1355 => x"54547281",
  1356 => x"2e9b3873",
  1357 => x"80c9dc0c",
  1358 => x"dfab3fdd",
  1359 => x"c33f80c1",
  1360 => x"e4528151",
  1361 => x"e4983fb0",
  1362 => x"0851879b",
  1363 => x"3f7280c9",
  1364 => x"dc0cdf91",
  1365 => x"3fdda93f",
  1366 => x"80c1e452",
  1367 => x"8151e3fe",
  1368 => x"3fb00851",
  1369 => x"87813f00",
  1370 => x"ff3900ff",
  1371 => x"39f53d0d",
  1372 => x"7e6080c9",
  1373 => x"dc08705b",
  1374 => x"585b5b75",
  1375 => x"80c23877",
  1376 => x"7a25a138",
  1377 => x"771b7033",
  1378 => x"7081ff06",
  1379 => x"58585975",
  1380 => x"8a2e9838",
  1381 => x"7681ff06",
  1382 => x"51dea93f",
  1383 => x"81185879",
  1384 => x"7824e138",
  1385 => x"79b00c8d",
  1386 => x"3d0d048d",
  1387 => x"51de953f",
  1388 => x"78337081",
  1389 => x"ff065257",
  1390 => x"de8a3f81",
  1391 => x"1858e039",
  1392 => x"79557a54",
  1393 => x"7d538552",
  1394 => x"8d3dfc05",
  1395 => x"51dcf23f",
  1396 => x"b0085686",
  1397 => x"8b3f7bb0",
  1398 => x"080c75b0",
  1399 => x"0c8d3d0d",
  1400 => x"04f63d0d",
  1401 => x"7d7f80c9",
  1402 => x"dc08705b",
  1403 => x"585a5a75",
  1404 => x"80c13877",
  1405 => x"7925b338",
  1406 => x"dda53fb0",
  1407 => x"0881ff06",
  1408 => x"708d3270",
  1409 => x"30709f2a",
  1410 => x"51515757",
  1411 => x"768a2e80",
  1412 => x"c3387580",
  1413 => x"2ebe3877",
  1414 => x"1a567676",
  1415 => x"347651dd",
  1416 => x"a33f8118",
  1417 => x"58787824",
  1418 => x"cf387756",
  1419 => x"75b00c8c",
  1420 => x"3d0d0478",
  1421 => x"5579547c",
  1422 => x"5384528c",
  1423 => x"3dfc0551",
  1424 => x"dbff3fb0",
  1425 => x"08568598",
  1426 => x"3f7ab008",
  1427 => x"0c75b00c",
  1428 => x"8c3d0d04",
  1429 => x"771a568a",
  1430 => x"76348118",
  1431 => x"588d51dc",
  1432 => x"e33f8a51",
  1433 => x"dcde3f77",
  1434 => x"56c239f9",
  1435 => x"3d0d7957",
  1436 => x"80c9dc08",
  1437 => x"802eac38",
  1438 => x"7651879e",
  1439 => x"3f7b567a",
  1440 => x"55b00881",
  1441 => x"05547653",
  1442 => x"8252893d",
  1443 => x"fc0551db",
  1444 => x"b03fb008",
  1445 => x"5784c93f",
  1446 => x"77b0080c",
  1447 => x"76b00c89",
  1448 => x"3d0d0484",
  1449 => x"bb3f850b",
  1450 => x"b0080cff",
  1451 => x"0bb00c89",
  1452 => x"3d0d04fb",
  1453 => x"3d0d80c9",
  1454 => x"dc087056",
  1455 => x"54738838",
  1456 => x"74b00c87",
  1457 => x"3d0d0477",
  1458 => x"53835287",
  1459 => x"3dfc0551",
  1460 => x"daef3fb0",
  1461 => x"08548488",
  1462 => x"3f75b008",
  1463 => x"0c73b00c",
  1464 => x"873d0d04",
  1465 => x"ff0bb00c",
  1466 => x"04fb3d0d",
  1467 => x"775580c9",
  1468 => x"dc08802e",
  1469 => x"a8387451",
  1470 => x"86a03fb0",
  1471 => x"08810554",
  1472 => x"74538752",
  1473 => x"873dfc05",
  1474 => x"51dab63f",
  1475 => x"b0085583",
  1476 => x"cf3f75b0",
  1477 => x"080c74b0",
  1478 => x"0c873d0d",
  1479 => x"0483c13f",
  1480 => x"850bb008",
  1481 => x"0cff0bb0",
  1482 => x"0c873d0d",
  1483 => x"04fa3d0d",
  1484 => x"80c9dc08",
  1485 => x"802ea238",
  1486 => x"7a557954",
  1487 => x"78538652",
  1488 => x"883dfc05",
  1489 => x"51d9fa3f",
  1490 => x"b0085683",
  1491 => x"933f76b0",
  1492 => x"080c75b0",
  1493 => x"0c883d0d",
  1494 => x"0483853f",
  1495 => x"9d0bb008",
  1496 => x"0cff0bb0",
  1497 => x"0c883d0d",
  1498 => x"04fb3d0d",
  1499 => x"77795656",
  1500 => x"80705454",
  1501 => x"7375259f",
  1502 => x"38741010",
  1503 => x"10f80552",
  1504 => x"72167033",
  1505 => x"70742b76",
  1506 => x"078116f8",
  1507 => x"16565656",
  1508 => x"51517473",
  1509 => x"24ea3873",
  1510 => x"b00c873d",
  1511 => x"0d04fc3d",
  1512 => x"0d767855",
  1513 => x"55bc5380",
  1514 => x"52735183",
  1515 => x"de3f8452",
  1516 => x"7451ffb5",
  1517 => x"3fb00874",
  1518 => x"23845284",
  1519 => x"1551ffa9",
  1520 => x"3fb00882",
  1521 => x"15238452",
  1522 => x"881551ff",
  1523 => x"9c3fb008",
  1524 => x"84150c84",
  1525 => x"528c1551",
  1526 => x"ff8f3fb0",
  1527 => x"08881523",
  1528 => x"84529015",
  1529 => x"51ff823f",
  1530 => x"b0088a15",
  1531 => x"23845294",
  1532 => x"1551fef5",
  1533 => x"3fb0088c",
  1534 => x"15238452",
  1535 => x"981551fe",
  1536 => x"e83fb008",
  1537 => x"8e152388",
  1538 => x"529c1551",
  1539 => x"fedb3fb0",
  1540 => x"0890150c",
  1541 => x"863d0d04",
  1542 => x"e93d0d6a",
  1543 => x"80c9dc08",
  1544 => x"57577593",
  1545 => x"3880c080",
  1546 => x"0b84180c",
  1547 => x"75ac180c",
  1548 => x"75b00c99",
  1549 => x"3d0d0489",
  1550 => x"3d70556a",
  1551 => x"54558a52",
  1552 => x"993dffbc",
  1553 => x"0551d7f9",
  1554 => x"3fb00877",
  1555 => x"53755256",
  1556 => x"fecc3f81",
  1557 => x"8b3f77b0",
  1558 => x"080c75b0",
  1559 => x"0c993d0d",
  1560 => x"04e93d0d",
  1561 => x"695780c9",
  1562 => x"dc08802e",
  1563 => x"b5387651",
  1564 => x"83a83f89",
  1565 => x"3d7056b0",
  1566 => x"08810555",
  1567 => x"7754568f",
  1568 => x"52993dff",
  1569 => x"bc0551d7",
  1570 => x"b83fb008",
  1571 => x"6b537652",
  1572 => x"57fe8b3f",
  1573 => x"80ca3f77",
  1574 => x"b0080c76",
  1575 => x"b00c993d",
  1576 => x"0d04bd3f",
  1577 => x"850bb008",
  1578 => x"0cff0bb0",
  1579 => x"0c993d0d",
  1580 => x"04fc3d0d",
  1581 => x"815480c9",
  1582 => x"dc088838",
  1583 => x"73b00c86",
  1584 => x"3d0d0476",
  1585 => x"5397b952",
  1586 => x"863dfc05",
  1587 => x"51d6f23f",
  1588 => x"b008548c",
  1589 => x"3f74b008",
  1590 => x"0c73b00c",
  1591 => x"863d0d04",
  1592 => x"80c1e808",
  1593 => x"b00c04f7",
  1594 => x"3d0d7b80",
  1595 => x"c1e80882",
  1596 => x"c811085a",
  1597 => x"545a7780",
  1598 => x"2e80da38",
  1599 => x"81881884",
  1600 => x"1908ff05",
  1601 => x"81712b59",
  1602 => x"55598074",
  1603 => x"2480ea38",
  1604 => x"807424b5",
  1605 => x"3873822b",
  1606 => x"78118805",
  1607 => x"56568180",
  1608 => x"19087706",
  1609 => x"5372802e",
  1610 => x"b6387816",
  1611 => x"70085353",
  1612 => x"79517408",
  1613 => x"53722dff",
  1614 => x"14fc17fc",
  1615 => x"1779812c",
  1616 => x"5a575754",
  1617 => x"738025d6",
  1618 => x"38770858",
  1619 => x"77ffad38",
  1620 => x"80c1e808",
  1621 => x"53bc1308",
  1622 => x"a5387951",
  1623 => x"f8893f74",
  1624 => x"0853722d",
  1625 => x"ff14fc17",
  1626 => x"fc177981",
  1627 => x"2c5a5757",
  1628 => x"54738025",
  1629 => x"ffa838d1",
  1630 => x"398057ff",
  1631 => x"93397251",
  1632 => x"bc130853",
  1633 => x"722d7951",
  1634 => x"f7dd3ffc",
  1635 => x"3d0d7679",
  1636 => x"71028c05",
  1637 => x"9f053357",
  1638 => x"55535583",
  1639 => x"72278a38",
  1640 => x"74830651",
  1641 => x"70802ea2",
  1642 => x"38ff1252",
  1643 => x"71ff2e93",
  1644 => x"38737370",
  1645 => x"81055534",
  1646 => x"ff125271",
  1647 => x"ff2e0981",
  1648 => x"06ef3874",
  1649 => x"b00c863d",
  1650 => x"0d047474",
  1651 => x"882b7507",
  1652 => x"7071902b",
  1653 => x"07515451",
  1654 => x"8f7227a5",
  1655 => x"38727170",
  1656 => x"8405530c",
  1657 => x"72717084",
  1658 => x"05530c72",
  1659 => x"71708405",
  1660 => x"530c7271",
  1661 => x"70840553",
  1662 => x"0cf01252",
  1663 => x"718f26dd",
  1664 => x"38837227",
  1665 => x"90387271",
  1666 => x"70840553",
  1667 => x"0cfc1252",
  1668 => x"718326f2",
  1669 => x"387053ff",
  1670 => x"9039fd3d",
  1671 => x"0d757071",
  1672 => x"83065355",
  1673 => x"5270b838",
  1674 => x"71700870",
  1675 => x"09f7fbfd",
  1676 => x"ff120670",
  1677 => x"f8848281",
  1678 => x"80065151",
  1679 => x"5253709d",
  1680 => x"38841370",
  1681 => x"087009f7",
  1682 => x"fbfdff12",
  1683 => x"0670f884",
  1684 => x"82818006",
  1685 => x"51515253",
  1686 => x"70802ee5",
  1687 => x"38725271",
  1688 => x"33517080",
  1689 => x"2e8a3881",
  1690 => x"12703352",
  1691 => x"5270f838",
  1692 => x"717431b0",
  1693 => x"0c853d0d",
  1694 => x"04ff3d0d",
  1695 => x"80c8ec0b",
  1696 => x"fc057008",
  1697 => x"525270ff",
  1698 => x"2e913870",
  1699 => x"2dfc1270",
  1700 => x"08525270",
  1701 => x"ff2e0981",
  1702 => x"06f13883",
  1703 => x"3d0d0404",
  1704 => x"d68b3f04",
  1705 => x"00ffffff",
  1706 => x"ff00ffff",
  1707 => x"ffff00ff",
  1708 => x"ffffff00",
  1709 => x"00000040",
  1710 => x"44485259",
  1711 => x"53544f4e",
  1712 => x"45205052",
  1713 => x"4f475241",
  1714 => x"4d2c2053",
  1715 => x"4f4d4520",
  1716 => x"53545249",
  1717 => x"4e470000",
  1718 => x"44485259",
  1719 => x"53544f4e",
  1720 => x"45205052",
  1721 => x"4f475241",
  1722 => x"4d2c2031",
  1723 => x"27535420",
  1724 => x"53545249",
  1725 => x"4e470000",
  1726 => x"44687279",
  1727 => x"73746f6e",
  1728 => x"65204265",
  1729 => x"6e63686d",
  1730 => x"61726b2c",
  1731 => x"20566572",
  1732 => x"73696f6e",
  1733 => x"20322e31",
  1734 => x"20284c61",
  1735 => x"6e677561",
  1736 => x"67653a20",
  1737 => x"43290a00",
  1738 => x"50726f67",
  1739 => x"72616d20",
  1740 => x"636f6d70",
  1741 => x"696c6564",
  1742 => x"20776974",
  1743 => x"68202772",
  1744 => x"65676973",
  1745 => x"74657227",
  1746 => x"20617474",
  1747 => x"72696275",
  1748 => x"74650a00",
  1749 => x"45786563",
  1750 => x"7574696f",
  1751 => x"6e207374",
  1752 => x"61727473",
  1753 => x"2c202564",
  1754 => x"2072756e",
  1755 => x"73207468",
  1756 => x"726f7567",
  1757 => x"68204468",
  1758 => x"72797374",
  1759 => x"6f6e650a",
  1760 => x"00000000",
  1761 => x"44485259",
  1762 => x"53544f4e",
  1763 => x"45205052",
  1764 => x"4f475241",
  1765 => x"4d2c2032",
  1766 => x"274e4420",
  1767 => x"53545249",
  1768 => x"4e470000",
  1769 => x"45786563",
  1770 => x"7574696f",
  1771 => x"6e20656e",
  1772 => x"64730a00",
  1773 => x"46696e61",
  1774 => x"6c207661",
  1775 => x"6c756573",
  1776 => x"206f6620",
  1777 => x"74686520",
  1778 => x"76617269",
  1779 => x"61626c65",
  1780 => x"73207573",
  1781 => x"65642069",
  1782 => x"6e207468",
  1783 => x"65206265",
  1784 => x"6e63686d",
  1785 => x"61726b3a",
  1786 => x"0a000000",
  1787 => x"496e745f",
  1788 => x"476c6f62",
  1789 => x"3a202020",
  1790 => x"20202020",
  1791 => x"20202020",
  1792 => x"2025640a",
  1793 => x"00000000",
  1794 => x"20202020",
  1795 => x"20202020",
  1796 => x"73686f75",
  1797 => x"6c642062",
  1798 => x"653a2020",
  1799 => x"2025640a",
  1800 => x"00000000",
  1801 => x"426f6f6c",
  1802 => x"5f476c6f",
  1803 => x"623a2020",
  1804 => x"20202020",
  1805 => x"20202020",
  1806 => x"2025640a",
  1807 => x"00000000",
  1808 => x"43685f31",
  1809 => x"5f476c6f",
  1810 => x"623a2020",
  1811 => x"20202020",
  1812 => x"20202020",
  1813 => x"2025630a",
  1814 => x"00000000",
  1815 => x"20202020",
  1816 => x"20202020",
  1817 => x"73686f75",
  1818 => x"6c642062",
  1819 => x"653a2020",
  1820 => x"2025630a",
  1821 => x"00000000",
  1822 => x"43685f32",
  1823 => x"5f476c6f",
  1824 => x"623a2020",
  1825 => x"20202020",
  1826 => x"20202020",
  1827 => x"2025630a",
  1828 => x"00000000",
  1829 => x"4172725f",
  1830 => x"315f476c",
  1831 => x"6f625b38",
  1832 => x"5d3a2020",
  1833 => x"20202020",
  1834 => x"2025640a",
  1835 => x"00000000",
  1836 => x"4172725f",
  1837 => x"325f476c",
  1838 => x"6f625b38",
  1839 => x"5d5b375d",
  1840 => x"3a202020",
  1841 => x"2025640a",
  1842 => x"00000000",
  1843 => x"20202020",
  1844 => x"20202020",
  1845 => x"73686f75",
  1846 => x"6c642062",
  1847 => x"653a2020",
  1848 => x"204e756d",
  1849 => x"6265725f",
  1850 => x"4f665f52",
  1851 => x"756e7320",
  1852 => x"2b203130",
  1853 => x"0a000000",
  1854 => x"5074725f",
  1855 => x"476c6f62",
  1856 => x"2d3e0a00",
  1857 => x"20205074",
  1858 => x"725f436f",
  1859 => x"6d703a20",
  1860 => x"20202020",
  1861 => x"20202020",
  1862 => x"2025640a",
  1863 => x"00000000",
  1864 => x"20202020",
  1865 => x"20202020",
  1866 => x"73686f75",
  1867 => x"6c642062",
  1868 => x"653a2020",
  1869 => x"2028696d",
  1870 => x"706c656d",
  1871 => x"656e7461",
  1872 => x"74696f6e",
  1873 => x"2d646570",
  1874 => x"656e6465",
  1875 => x"6e74290a",
  1876 => x"00000000",
  1877 => x"20204469",
  1878 => x"7363723a",
  1879 => x"20202020",
  1880 => x"20202020",
  1881 => x"20202020",
  1882 => x"2025640a",
  1883 => x"00000000",
  1884 => x"2020456e",
  1885 => x"756d5f43",
  1886 => x"6f6d703a",
  1887 => x"20202020",
  1888 => x"20202020",
  1889 => x"2025640a",
  1890 => x"00000000",
  1891 => x"2020496e",
  1892 => x"745f436f",
  1893 => x"6d703a20",
  1894 => x"20202020",
  1895 => x"20202020",
  1896 => x"2025640a",
  1897 => x"00000000",
  1898 => x"20205374",
  1899 => x"725f436f",
  1900 => x"6d703a20",
  1901 => x"20202020",
  1902 => x"20202020",
  1903 => x"2025730a",
  1904 => x"00000000",
  1905 => x"20202020",
  1906 => x"20202020",
  1907 => x"73686f75",
  1908 => x"6c642062",
  1909 => x"653a2020",
  1910 => x"20444852",
  1911 => x"5953544f",
  1912 => x"4e452050",
  1913 => x"524f4752",
  1914 => x"414d2c20",
  1915 => x"534f4d45",
  1916 => x"20535452",
  1917 => x"494e470a",
  1918 => x"00000000",
  1919 => x"4e657874",
  1920 => x"5f507472",
  1921 => x"5f476c6f",
  1922 => x"622d3e0a",
  1923 => x"00000000",
  1924 => x"20202020",
  1925 => x"20202020",
  1926 => x"73686f75",
  1927 => x"6c642062",
  1928 => x"653a2020",
  1929 => x"2028696d",
  1930 => x"706c656d",
  1931 => x"656e7461",
  1932 => x"74696f6e",
  1933 => x"2d646570",
  1934 => x"656e6465",
  1935 => x"6e74292c",
  1936 => x"2073616d",
  1937 => x"65206173",
  1938 => x"2061626f",
  1939 => x"76650a00",
  1940 => x"496e745f",
  1941 => x"315f4c6f",
  1942 => x"633a2020",
  1943 => x"20202020",
  1944 => x"20202020",
  1945 => x"2025640a",
  1946 => x"00000000",
  1947 => x"496e745f",
  1948 => x"325f4c6f",
  1949 => x"633a2020",
  1950 => x"20202020",
  1951 => x"20202020",
  1952 => x"2025640a",
  1953 => x"00000000",
  1954 => x"496e745f",
  1955 => x"335f4c6f",
  1956 => x"633a2020",
  1957 => x"20202020",
  1958 => x"20202020",
  1959 => x"2025640a",
  1960 => x"00000000",
  1961 => x"456e756d",
  1962 => x"5f4c6f63",
  1963 => x"3a202020",
  1964 => x"20202020",
  1965 => x"20202020",
  1966 => x"2025640a",
  1967 => x"00000000",
  1968 => x"5374725f",
  1969 => x"315f4c6f",
  1970 => x"633a2020",
  1971 => x"20202020",
  1972 => x"20202020",
  1973 => x"2025730a",
  1974 => x"00000000",
  1975 => x"20202020",
  1976 => x"20202020",
  1977 => x"73686f75",
  1978 => x"6c642062",
  1979 => x"653a2020",
  1980 => x"20444852",
  1981 => x"5953544f",
  1982 => x"4e452050",
  1983 => x"524f4752",
  1984 => x"414d2c20",
  1985 => x"31275354",
  1986 => x"20535452",
  1987 => x"494e470a",
  1988 => x"00000000",
  1989 => x"5374725f",
  1990 => x"325f4c6f",
  1991 => x"633a2020",
  1992 => x"20202020",
  1993 => x"20202020",
  1994 => x"2025730a",
  1995 => x"00000000",
  1996 => x"20202020",
  1997 => x"20202020",
  1998 => x"73686f75",
  1999 => x"6c642062",
  2000 => x"653a2020",
  2001 => x"20444852",
  2002 => x"5953544f",
  2003 => x"4e452050",
  2004 => x"524f4752",
  2005 => x"414d2c20",
  2006 => x"32274e44",
  2007 => x"20535452",
  2008 => x"494e470a",
  2009 => x"00000000",
  2010 => x"55736572",
  2011 => x"2074696d",
  2012 => x"653a2025",
  2013 => x"640a0000",
  2014 => x"4d696372",
  2015 => x"6f736563",
  2016 => x"6f6e6473",
  2017 => x"20666f72",
  2018 => x"206f6e65",
  2019 => x"2072756e",
  2020 => x"20746872",
  2021 => x"6f756768",
  2022 => x"20446872",
  2023 => x"7973746f",
  2024 => x"6e653a20",
  2025 => x"00000000",
  2026 => x"2564200a",
  2027 => x"00000000",
  2028 => x"44687279",
  2029 => x"73746f6e",
  2030 => x"65732070",
  2031 => x"65722053",
  2032 => x"65636f6e",
  2033 => x"643a2020",
  2034 => x"20202020",
  2035 => x"20202020",
  2036 => x"20202020",
  2037 => x"20202020",
  2038 => x"20202020",
  2039 => x"00000000",
  2040 => x"56415820",
  2041 => x"4d495053",
  2042 => x"20726174",
  2043 => x"696e6720",
  2044 => x"2a203130",
  2045 => x"3030203d",
  2046 => x"20256420",
  2047 => x"0a000000",
  2048 => x"50726f67",
  2049 => x"72616d20",
  2050 => x"636f6d70",
  2051 => x"696c6564",
  2052 => x"20776974",
  2053 => x"686f7574",
  2054 => x"20277265",
  2055 => x"67697374",
  2056 => x"65722720",
  2057 => x"61747472",
  2058 => x"69627574",
  2059 => x"650a0000",
  2060 => x"4d656173",
  2061 => x"75726564",
  2062 => x"2074696d",
  2063 => x"6520746f",
  2064 => x"6f20736d",
  2065 => x"616c6c20",
  2066 => x"746f206f",
  2067 => x"62746169",
  2068 => x"6e206d65",
  2069 => x"616e696e",
  2070 => x"6766756c",
  2071 => x"20726573",
  2072 => x"756c7473",
  2073 => x"0a000000",
  2074 => x"506c6561",
  2075 => x"73652069",
  2076 => x"6e637265",
  2077 => x"61736520",
  2078 => x"6e756d62",
  2079 => x"6572206f",
  2080 => x"66207275",
  2081 => x"6e730a00",
  2082 => x"44485259",
  2083 => x"53544f4e",
  2084 => x"45205052",
  2085 => x"4f475241",
  2086 => x"4d2c2033",
  2087 => x"27524420",
  2088 => x"53545249",
  2089 => x"4e470000",
  2090 => x"30313233",
  2091 => x"34353637",
  2092 => x"38394142",
  2093 => x"43444546",
  2094 => x"00000000",
  2095 => x"64756d6d",
  2096 => x"792e6578",
  2097 => x"65000000",
  2098 => x"43000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00002474",
  2103 => x"000061a8",
  2104 => x"00000000",
  2105 => x"000020bc",
  2106 => x"000020ec",
  2107 => x"00000000",
  2108 => x"00002354",
  2109 => x"000023b0",
  2110 => x"0000240c",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"000020c8",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000001",
  2150 => x"330eabcd",
  2151 => x"1234e66d",
  2152 => x"deec0005",
  2153 => x"000b0000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"00000000",
  2209 => x"00000000",
  2210 => x"00000000",
  2211 => x"00000000",
  2212 => x"00000000",
  2213 => x"00000000",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"00000000",
  2217 => x"00000000",
  2218 => x"00000000",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000000",
  2244 => x"00000000",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"00000000",
  2262 => x"00000000",
  2263 => x"00000000",
  2264 => x"00000000",
  2265 => x"00000000",
  2266 => x"00000000",
  2267 => x"00000000",
  2268 => x"00000000",
  2269 => x"00000000",
  2270 => x"00000000",
  2271 => x"00000000",
  2272 => x"00000000",
  2273 => x"00000000",
  2274 => x"00000000",
  2275 => x"00000000",
  2276 => x"00000000",
  2277 => x"00000000",
  2278 => x"00000000",
  2279 => x"00000000",
  2280 => x"00000000",
  2281 => x"00000000",
  2282 => x"00000000",
  2283 => x"00000000",
  2284 => x"00000000",
  2285 => x"00000000",
  2286 => x"00000000",
  2287 => x"00000000",
  2288 => x"00000000",
  2289 => x"00000000",
  2290 => x"00000000",
  2291 => x"00000000",
  2292 => x"00000000",
  2293 => x"00000000",
  2294 => x"00000000",
  2295 => x"00000000",
  2296 => x"00000000",
  2297 => x"00000000",
  2298 => x"00000000",
  2299 => x"00000000",
  2300 => x"00000000",
  2301 => x"00000000",
  2302 => x"00000000",
  2303 => x"00000000",
  2304 => x"00000000",
  2305 => x"00000000",
  2306 => x"00000000",
  2307 => x"00000000",
  2308 => x"00000000",
  2309 => x"00000000",
  2310 => x"00000000",
  2311 => x"00000000",
  2312 => x"00000000",
  2313 => x"00000000",
  2314 => x"00000000",
  2315 => x"00000000",
  2316 => x"00000000",
  2317 => x"00000000",
  2318 => x"00000000",
  2319 => x"00000000",
  2320 => x"00000000",
  2321 => x"00000000",
  2322 => x"00000000",
  2323 => x"00000000",
  2324 => x"00000000",
  2325 => x"00000000",
  2326 => x"00000000",
  2327 => x"00000000",
  2328 => x"00000000",
  2329 => x"00000000",
  2330 => x"ffffffff",
  2331 => x"00000000",
  2332 => x"ffffffff",
  2333 => x"00000000",
  2334 => x"00000000",
	others => x"00000000"
);

begin

mem_busy<=mem_readEnable; -- we're done on the cycle after we serve the read request

process (clk, areset)
begin
		if areset = '1' then
		elsif (clk'event and clk = '1') then
			if (mem_writeEnable = '1') then
				ram(to_integer(unsigned(mem_addr(maxAddrBit downto minAddrBit)))) := mem_write;
			end if;
		if (mem_readEnable = '1') then
			mem_read <= ram(to_integer(unsigned(mem_addr(maxAddrBit downto minAddrBit))));
		end if;
	end if;
end process;




end dram_arch;


-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"f2040000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"97a07383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040ba0",
    29 => x"8080fd0b",
    30 => x"a080888d",
    31 => x"040ba080",
    32 => x"80fd0402",
    33 => x"f4050d74",
    34 => x"767181ff",
    35 => x"06c80c53",
    36 => x"5383fff0",
    37 => x"9c088538",
    38 => x"71892b52",
    39 => x"71982ac8",
    40 => x"0c71902a",
    41 => x"7081ff06",
    42 => x"c80c5171",
    43 => x"882a7081",
    44 => x"ff06c80c",
    45 => x"517181ff",
    46 => x"06c80c72",
    47 => x"902a7081",
    48 => x"ff06c80c",
    49 => x"51c80870",
    50 => x"81ff0651",
    51 => x"5182b8bf",
    52 => x"527081ff",
    53 => x"2e098106",
    54 => x"943881ff",
    55 => x"0bc80cc8",
    56 => x"087081ff",
    57 => x"06ff1454",
    58 => x"515171e5",
    59 => x"387083ff",
    60 => x"e0800c02",
    61 => x"8c050d04",
    62 => x"02fc050d",
    63 => x"81c75181",
    64 => x"ff0bc80c",
    65 => x"ff115170",
    66 => x"8025f438",
    67 => x"0284050d",
    68 => x"0402f005",
    69 => x"0da08081",
    70 => x"f82d819c",
    71 => x"9f538052",
    72 => x"87fc80f7",
    73 => x"51a08081",
    74 => x"832d83ff",
    75 => x"e0800854",
    76 => x"83ffe080",
    77 => x"08812e09",
    78 => x"8106ab38",
    79 => x"81ff0bc8",
    80 => x"0c820a52",
    81 => x"849c80e9",
    82 => x"51a08081",
    83 => x"832d83ff",
    84 => x"e080088d",
    85 => x"3881ff0b",
    86 => x"c80c7353",
    87 => x"a08082ed",
    88 => x"04a08081",
    89 => x"f82dff13",
    90 => x"5372ffb2",
    91 => x"387283ff",
    92 => x"e0800c02",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"81ff0bc8",
    96 => x"0c935380",
    97 => x"5287fc80",
    98 => x"c151a080",
    99 => x"81832d83",
   100 => x"ffe08008",
   101 => x"8d3881ff",
   102 => x"0bc80c81",
   103 => x"53a08083",
   104 => x"ad04a080",
   105 => x"81f82dff",
   106 => x"135372d7",
   107 => x"387283ff",
   108 => x"e0800c02",
   109 => x"8c050d04",
   110 => x"02f0050d",
   111 => x"a08081f8",
   112 => x"2d83aa52",
   113 => x"849c80c8",
   114 => x"51a08081",
   115 => x"832d83ff",
   116 => x"e0800881",
   117 => x"2e098106",
   118 => x"9038cc08",
   119 => x"7083ffff",
   120 => x"06515372",
   121 => x"83aa2e99",
   122 => x"38a08082",
   123 => x"f82da080",
   124 => x"83fa0481",
   125 => x"54a08084",
   126 => x"db048054",
   127 => x"a08084db",
   128 => x"0481ff0b",
   129 => x"c80cb153",
   130 => x"a0808291",
   131 => x"2d83ffe0",
   132 => x"8008802e",
   133 => x"b7388052",
   134 => x"87fc80fa",
   135 => x"51a08081",
   136 => x"832d83ff",
   137 => x"e08008a4",
   138 => x"3881ff0b",
   139 => x"c80cc808",
   140 => x"cc087186",
   141 => x"2a708106",
   142 => x"83ffe080",
   143 => x"08535152",
   144 => x"55537280",
   145 => x"2e9538a0",
   146 => x"8083f304",
   147 => x"72822eff",
   148 => x"a938ff13",
   149 => x"5372ffb0",
   150 => x"38725473",
   151 => x"83ffe080",
   152 => x"0c029005",
   153 => x"0d0402f4",
   154 => x"050d810b",
   155 => x"83fff09c",
   156 => x"0cc40870",
   157 => x"8f2a7081",
   158 => x"06515153",
   159 => x"72f33872",
   160 => x"c40ca080",
   161 => x"81f82dc4",
   162 => x"08708f2a",
   163 => x"70810651",
   164 => x"515372f3",
   165 => x"38810bc4",
   166 => x"0c875380",
   167 => x"5284d480",
   168 => x"c051a080",
   169 => x"81832d83",
   170 => x"ffe08008",
   171 => x"812e9638",
   172 => x"72822e09",
   173 => x"81068838",
   174 => x"8053a080",
   175 => x"85fd04ff",
   176 => x"135372d7",
   177 => x"38a08083",
   178 => x"b82d83ff",
   179 => x"e0800883",
   180 => x"fff09c0c",
   181 => x"815287fc",
   182 => x"80d051a0",
   183 => x"8081832d",
   184 => x"81ff0bc8",
   185 => x"0cc40870",
   186 => x"8f2a7081",
   187 => x"06515153",
   188 => x"72f33872",
   189 => x"c40c81ff",
   190 => x"0bc80c81",
   191 => x"537283ff",
   192 => x"e0800c02",
   193 => x"8c050d04",
   194 => x"800b83ff",
   195 => x"e0800c04",
   196 => x"02e8050d",
   197 => x"78558056",
   198 => x"c408708f",
   199 => x"2a708106",
   200 => x"51515372",
   201 => x"f3388281",
   202 => x"0bc40c81",
   203 => x"ff0bc80c",
   204 => x"775287fc",
   205 => x"80d151a0",
   206 => x"8081832d",
   207 => x"83ffe080",
   208 => x"0880d238",
   209 => x"80dbc6df",
   210 => x"5481ff0b",
   211 => x"c80cc808",
   212 => x"7081ff06",
   213 => x"51537281",
   214 => x"fe2e0981",
   215 => x"069b3880",
   216 => x"ff54cc08",
   217 => x"75708405",
   218 => x"570cff14",
   219 => x"54738025",
   220 => x"f1388156",
   221 => x"a08086ff",
   222 => x"04ff1454",
   223 => x"73cb3881",
   224 => x"ff0bc80c",
   225 => x"c408708f",
   226 => x"2a708106",
   227 => x"51515372",
   228 => x"f33872c4",
   229 => x"0c7583ff",
   230 => x"e0800c02",
   231 => x"98050d04",
   232 => x"02f4050d",
   233 => x"7470882a",
   234 => x"83fe8006",
   235 => x"7072982a",
   236 => x"0772882b",
   237 => x"87fc8080",
   238 => x"0673982b",
   239 => x"81f00a06",
   240 => x"71730707",
   241 => x"83ffe080",
   242 => x"0c565153",
   243 => x"51028c05",
   244 => x"0d0402f4",
   245 => x"050d0292",
   246 => x"05a08080",
   247 => x"9f2d7088",
   248 => x"2a71882b",
   249 => x"077083ff",
   250 => x"ff0683ff",
   251 => x"e0800c52",
   252 => x"52028c05",
   253 => x"0d0402f8",
   254 => x"050d7370",
   255 => x"902b7190",
   256 => x"2a0783ff",
   257 => x"e0800c52",
   258 => x"0288050d",
   259 => x"0402ec05",
   260 => x"0d88bd0b",
   261 => x"ff880c80",
   262 => x"0b870a0c",
   263 => x"f80883ff",
   264 => x"f0900cfc",
   265 => x"0883fff0",
   266 => x"940c84ea",
   267 => x"cda8800b",
   268 => x"83fff098",
   269 => x"0ca08084",
   270 => x"e62d83ff",
   271 => x"e0800880",
   272 => x"2e81d138",
   273 => x"a0808ae8",
   274 => x"2d83ffe0",
   275 => x"905283ff",
   276 => x"f09051a0",
   277 => x"8095ed2d",
   278 => x"83ffe080",
   279 => x"08802e81",
   280 => x"b33883ff",
   281 => x"e0905480",
   282 => x"55737081",
   283 => x"0555a080",
   284 => x"80b42d53",
   285 => x"72a02e80",
   286 => x"de3872a3",
   287 => x"2e80fd38",
   288 => x"7280c72e",
   289 => x"0981068b",
   290 => x"38a08080",
   291 => x"882da080",
   292 => x"89b30472",
   293 => x"8a2e0981",
   294 => x"068b38a0",
   295 => x"8080902d",
   296 => x"a08089b3",
   297 => x"047280cc",
   298 => x"2e098106",
   299 => x"863883ff",
   300 => x"e0905472",
   301 => x"81df06f0",
   302 => x"057081ff",
   303 => x"065153b8",
   304 => x"73278938",
   305 => x"ef137081",
   306 => x"ff065153",
   307 => x"74842b73",
   308 => x"0755a080",
   309 => x"88e90472",
   310 => x"a32ea138",
   311 => x"73708105",
   312 => x"55a08080",
   313 => x"b42d5372",
   314 => x"a02ef138",
   315 => x"ff147553",
   316 => x"705254a0",
   317 => x"8095ed2d",
   318 => x"74870a0c",
   319 => x"73708105",
   320 => x"55a08080",
   321 => x"b42d5372",
   322 => x"8a2e0981",
   323 => x"06ee38a0",
   324 => x"8088e704",
   325 => x"800b83ff",
   326 => x"e0800c02",
   327 => x"94050d04",
   328 => x"02e8050d",
   329 => x"77797b58",
   330 => x"55558053",
   331 => x"727625ab",
   332 => x"38747081",
   333 => x"0556a080",
   334 => x"80b42d74",
   335 => x"70810556",
   336 => x"a08080b4",
   337 => x"2d525271",
   338 => x"712e8838",
   339 => x"8151a080",
   340 => x"8add0481",
   341 => x"1353a080",
   342 => x"8aac0480",
   343 => x"517083ff",
   344 => x"e0800c02",
   345 => x"98050d04",
   346 => x"02d8050d",
   347 => x"ff0b83ff",
   348 => x"f4c80c80",
   349 => x"0b83fff4",
   350 => x"dc0c83ff",
   351 => x"f0b45280",
   352 => x"51a08086",
   353 => x"902d83ff",
   354 => x"e0800855",
   355 => x"83ffe080",
   356 => x"08802e86",
   357 => x"d3388056",
   358 => x"810b83ff",
   359 => x"f0a80c88",
   360 => x"53a08097",
   361 => x"b05283ff",
   362 => x"f0ea51a0",
   363 => x"808aa02d",
   364 => x"83ffe080",
   365 => x"08762e09",
   366 => x"81068b38",
   367 => x"83ffe080",
   368 => x"0883fff0",
   369 => x"a80c8853",
   370 => x"a08097bc",
   371 => x"5283fff1",
   372 => x"8651a080",
   373 => x"8aa02d83",
   374 => x"ffe08008",
   375 => x"8b3883ff",
   376 => x"e0800883",
   377 => x"fff0a80c",
   378 => x"83fff0a8",
   379 => x"08802e81",
   380 => x"9c3883ff",
   381 => x"f3fa0ba0",
   382 => x"8080b42d",
   383 => x"83fff3fb",
   384 => x"0ba08080",
   385 => x"b42d7198",
   386 => x"2b71902b",
   387 => x"0783fff3",
   388 => x"fc0ba080",
   389 => x"80b42d70",
   390 => x"882b7207",
   391 => x"83fff3fd",
   392 => x"0ba08080",
   393 => x"b42d7107",
   394 => x"83fff4b2",
   395 => x"0ba08080",
   396 => x"b42d83ff",
   397 => x"f4b30ba0",
   398 => x"8080b42d",
   399 => x"71882b07",
   400 => x"535f5452",
   401 => x"5a565755",
   402 => x"7381abaa",
   403 => x"2e098106",
   404 => x"93387551",
   405 => x"a08087a0",
   406 => x"2d83ffe0",
   407 => x"800856a0",
   408 => x"808cf104",
   409 => x"80557382",
   410 => x"d4d52e09",
   411 => x"810684f8",
   412 => x"3883fff0",
   413 => x"b4527551",
   414 => x"a0808690",
   415 => x"2d83ffe0",
   416 => x"80085583",
   417 => x"ffe08008",
   418 => x"802e84dc",
   419 => x"388853a0",
   420 => x"8097bc52",
   421 => x"83fff186",
   422 => x"51a0808a",
   423 => x"a02d83ff",
   424 => x"e080088d",
   425 => x"38810b83",
   426 => x"fff4dc0c",
   427 => x"a0808dd1",
   428 => x"048853a0",
   429 => x"8097b052",
   430 => x"83fff0ea",
   431 => x"51a0808a",
   432 => x"a02d8055",
   433 => x"83ffe080",
   434 => x"08752e09",
   435 => x"81068498",
   436 => x"3883fff4",
   437 => x"b20ba080",
   438 => x"80b42d54",
   439 => x"7380d52e",
   440 => x"09810680",
   441 => x"db3883ff",
   442 => x"f4b30ba0",
   443 => x"8080b42d",
   444 => x"547381aa",
   445 => x"2e098106",
   446 => x"80c63880",
   447 => x"0b83fff0",
   448 => x"b40ba080",
   449 => x"80b42d56",
   450 => x"547481e9",
   451 => x"2e833881",
   452 => x"547481eb",
   453 => x"2e8c3880",
   454 => x"5573752e",
   455 => x"09810683",
   456 => x"c73883ff",
   457 => x"f0bf0ba0",
   458 => x"8080b42d",
   459 => x"55749138",
   460 => x"83fff0c0",
   461 => x"0ba08080",
   462 => x"b42d5473",
   463 => x"822e8838",
   464 => x"8055a080",
   465 => x"91e80483",
   466 => x"fff0c10b",
   467 => x"a08080b4",
   468 => x"2d7083ff",
   469 => x"f4e40cff",
   470 => x"0583fff4",
   471 => x"d80c83ff",
   472 => x"f0c20ba0",
   473 => x"8080b42d",
   474 => x"83fff0c3",
   475 => x"0ba08080",
   476 => x"b42d5876",
   477 => x"05778280",
   478 => x"29057083",
   479 => x"fff4cc0c",
   480 => x"83fff0c4",
   481 => x"0ba08080",
   482 => x"b42d7083",
   483 => x"fff4c40c",
   484 => x"83fff4dc",
   485 => x"08595758",
   486 => x"76802e81",
   487 => x"df388853",
   488 => x"a08097bc",
   489 => x"5283fff1",
   490 => x"8651a080",
   491 => x"8aa02d83",
   492 => x"ffe08008",
   493 => x"82b23883",
   494 => x"fff4e408",
   495 => x"70842b83",
   496 => x"fff4b40c",
   497 => x"7083fff4",
   498 => x"e00c83ff",
   499 => x"f0d90ba0",
   500 => x"8080b42d",
   501 => x"83fff0d8",
   502 => x"0ba08080",
   503 => x"b42d7182",
   504 => x"80290583",
   505 => x"fff0da0b",
   506 => x"a08080b4",
   507 => x"2d708480",
   508 => x"80291283",
   509 => x"fff0db0b",
   510 => x"a08080b4",
   511 => x"2d708180",
   512 => x"0a291270",
   513 => x"83fff0ac",
   514 => x"0c83fff4",
   515 => x"c4087129",
   516 => x"83fff4cc",
   517 => x"08057083",
   518 => x"fff4ec0c",
   519 => x"83fff0e1",
   520 => x"0ba08080",
   521 => x"b42d83ff",
   522 => x"f0e00ba0",
   523 => x"8080b42d",
   524 => x"71828029",
   525 => x"0583fff0",
   526 => x"e20ba080",
   527 => x"80b42d70",
   528 => x"84808029",
   529 => x"1283fff0",
   530 => x"e30ba080",
   531 => x"80b42d70",
   532 => x"982b81f0",
   533 => x"0a067205",
   534 => x"7083fff0",
   535 => x"b00cfe11",
   536 => x"7e297705",
   537 => x"83fff4d4",
   538 => x"0c525952",
   539 => x"43545e51",
   540 => x"5259525d",
   541 => x"575957a0",
   542 => x"8091e604",
   543 => x"83fff0c6",
   544 => x"0ba08080",
   545 => x"b42d83ff",
   546 => x"f0c50ba0",
   547 => x"8080b42d",
   548 => x"71828029",
   549 => x"057083ff",
   550 => x"f4b40c70",
   551 => x"a02983ff",
   552 => x"0570892a",
   553 => x"7083fff4",
   554 => x"e00c83ff",
   555 => x"f0cb0ba0",
   556 => x"8080b42d",
   557 => x"83fff0ca",
   558 => x"0ba08080",
   559 => x"b42d7182",
   560 => x"80290570",
   561 => x"83fff0ac",
   562 => x"0c7b7129",
   563 => x"1e7083ff",
   564 => x"f4d40c7d",
   565 => x"83fff0b0",
   566 => x"0c730583",
   567 => x"fff4ec0c",
   568 => x"555e5151",
   569 => x"55558155",
   570 => x"7483ffe0",
   571 => x"800c02a8",
   572 => x"050d0402",
   573 => x"ec050d76",
   574 => x"70872c71",
   575 => x"80ff0657",
   576 => x"555383ff",
   577 => x"f4dc088a",
   578 => x"3872882c",
   579 => x"7381ff06",
   580 => x"56547383",
   581 => x"fff4c808",
   582 => x"2ea83883",
   583 => x"fff0b452",
   584 => x"83fff4cc",
   585 => x"081451a0",
   586 => x"8086902d",
   587 => x"83ffe080",
   588 => x"085383ff",
   589 => x"e0800880",
   590 => x"2e80cb38",
   591 => x"7383fff4",
   592 => x"c80c83ff",
   593 => x"f4dc0880",
   594 => x"2ea03874",
   595 => x"842983ff",
   596 => x"f0b40570",
   597 => x"085253a0",
   598 => x"8087a02d",
   599 => x"83ffe080",
   600 => x"08f00a06",
   601 => x"55a08093",
   602 => x"84047410",
   603 => x"83fff0b4",
   604 => x"0570a080",
   605 => x"809f2d52",
   606 => x"53a08087",
   607 => x"d22d83ff",
   608 => x"e0800855",
   609 => x"74537283",
   610 => x"ffe0800c",
   611 => x"0294050d",
   612 => x"0402cc05",
   613 => x"0d7e605e",
   614 => x"5b8056ff",
   615 => x"0b83fff4",
   616 => x"c80c83ff",
   617 => x"f0b00883",
   618 => x"fff4d408",
   619 => x"565a83ff",
   620 => x"f4dc0876",
   621 => x"2e8e3883",
   622 => x"fff4e408",
   623 => x"842b58a0",
   624 => x"8093cc04",
   625 => x"83fff4e0",
   626 => x"08842b58",
   627 => x"80597878",
   628 => x"2781c938",
   629 => x"788f06a0",
   630 => x"17575473",
   631 => x"953883ff",
   632 => x"f0b45274",
   633 => x"51811555",
   634 => x"a0808690",
   635 => x"2d83fff0",
   636 => x"b4568076",
   637 => x"a08080b4",
   638 => x"2d555773",
   639 => x"772e8338",
   640 => x"81577381",
   641 => x"e52e818c",
   642 => x"38817078",
   643 => x"06555c73",
   644 => x"802e8180",
   645 => x"388b16a0",
   646 => x"8080b42d",
   647 => x"98065776",
   648 => x"80f2388b",
   649 => x"537c5275",
   650 => x"51a0808a",
   651 => x"a02d83ff",
   652 => x"e0800880",
   653 => x"df389c16",
   654 => x"0851a080",
   655 => x"87a02d83",
   656 => x"ffe08008",
   657 => x"841c0c9a",
   658 => x"16a08080",
   659 => x"9f2d51a0",
   660 => x"8087d22d",
   661 => x"83ffe080",
   662 => x"0883ffe0",
   663 => x"80085555",
   664 => x"83fff4dc",
   665 => x"08802e9e",
   666 => x"389416a0",
   667 => x"80809f2d",
   668 => x"51a08087",
   669 => x"d22d83ff",
   670 => x"e0800890",
   671 => x"2b83fff0",
   672 => x"0a067016",
   673 => x"51547388",
   674 => x"1c0c767b",
   675 => x"0c7b54a0",
   676 => x"8095e204",
   677 => x"811959a0",
   678 => x"8093ce04",
   679 => x"83fff4dc",
   680 => x"08802ebc",
   681 => x"387951a0",
   682 => x"8091f32d",
   683 => x"83ffe080",
   684 => x"0883ffe0",
   685 => x"800880ff",
   686 => x"fffff806",
   687 => x"555a7380",
   688 => x"fffffff8",
   689 => x"2e9a3883",
   690 => x"ffe08008",
   691 => x"fe0583ff",
   692 => x"f4e40829",
   693 => x"83fff4ec",
   694 => x"080555a0",
   695 => x"8093cc04",
   696 => x"80547383",
   697 => x"ffe0800c",
   698 => x"02b4050d",
   699 => x"0402e405",
   700 => x"0d797953",
   701 => x"83fff4b8",
   702 => x"5255a080",
   703 => x"93912d83",
   704 => x"ffe08008",
   705 => x"81ff0670",
   706 => x"55537280",
   707 => x"2e818538",
   708 => x"83fff4bc",
   709 => x"0883ff05",
   710 => x"892a5780",
   711 => x"70555675",
   712 => x"772580ee",
   713 => x"3883fff4",
   714 => x"c008fe05",
   715 => x"83fff4e4",
   716 => x"082983ff",
   717 => x"f4ec0811",
   718 => x"7583fff4",
   719 => x"d8080605",
   720 => x"76545253",
   721 => x"a0808690",
   722 => x"2d83ffe0",
   723 => x"8008802e",
   724 => x"b6388114",
   725 => x"7083fff4",
   726 => x"d8080654",
   727 => x"54729638",
   728 => x"83fff4c0",
   729 => x"0851a080",
   730 => x"91f32d83",
   731 => x"ffe08008",
   732 => x"83fff4c0",
   733 => x"0c848015",
   734 => x"81175755",
   735 => x"767624ff",
   736 => x"a438a080",
   737 => x"97920483",
   738 => x"ffe08008",
   739 => x"54a08097",
   740 => x"94048154",
   741 => x"7383ffe0",
   742 => x"800c029c",
   743 => x"050d0400",
   744 => x"00ffffff",
   745 => x"ff00ffff",
   746 => x"ffff00ff",
   747 => x"ffffff00",
   748 => x"46415431",
   749 => x"36202020",
   750 => x"00000000",
   751 => x"46415433",
   752 => x"32202020",
   753 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;


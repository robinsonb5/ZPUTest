-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dhrystone_rom is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end dhrystone_rom;

architecture arch of dhrystone_rom is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"80700b0b",
     2 => x"0bbff80c",
     3 => x"3a0b0b0b",
     4 => x"a8ca0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"8f040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bb3",
   162 => x"cc738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f7040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"df040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bbff40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"83df3fab",
   257 => x"9a3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104b0",
   280 => x"08b408b8",
   281 => x"087575a2",
   282 => x"f02d5050",
   283 => x"b00856b8",
   284 => x"0cb40cb0",
   285 => x"0c5104b0",
   286 => x"08b408b8",
   287 => x"087575a1",
   288 => x"be2d5050",
   289 => x"b00856b8",
   290 => x"0cb40cb0",
   291 => x"0c5104b0",
   292 => x"08b408b8",
   293 => x"08a9902d",
   294 => x"b80cb40c",
   295 => x"b00c04fe",
   296 => x"3d0d0b0b",
   297 => x"80c7a408",
   298 => x"53841308",
   299 => x"70882a70",
   300 => x"81065152",
   301 => x"5270802e",
   302 => x"f0387181",
   303 => x"ff06b00c",
   304 => x"843d0d04",
   305 => x"ff3d0d0b",
   306 => x"0b80c7a4",
   307 => x"08527108",
   308 => x"70882a81",
   309 => x"32708106",
   310 => x"51515170",
   311 => x"f1387372",
   312 => x"0c833d0d",
   313 => x"04bff408",
   314 => x"802ea338",
   315 => x"bff80882",
   316 => x"2ebd3883",
   317 => x"80800b0b",
   318 => x"0b80c7a4",
   319 => x"0c82a080",
   320 => x"0b80c7a8",
   321 => x"0c829080",
   322 => x"0b80c7ac",
   323 => x"0c04f880",
   324 => x"8080a40b",
   325 => x"0b0b80c7",
   326 => x"a40cf880",
   327 => x"8082800b",
   328 => x"80c7a80c",
   329 => x"f8808084",
   330 => x"800b80c7",
   331 => x"ac0c0480",
   332 => x"c0a8808c",
   333 => x"0b0b0b80",
   334 => x"c7a40c80",
   335 => x"c0a88094",
   336 => x"0b80c7a8",
   337 => x"0cb3dc0b",
   338 => x"80c7ac0c",
   339 => x"04f23d0d",
   340 => x"6080c7a8",
   341 => x"08565d82",
   342 => x"750c8059",
   343 => x"805a800b",
   344 => x"8f3d5d5b",
   345 => x"7a101015",
   346 => x"70087108",
   347 => x"719f2c7e",
   348 => x"852b5855",
   349 => x"557d5359",
   350 => x"5794cd3f",
   351 => x"7d7f7a72",
   352 => x"077c7207",
   353 => x"71716081",
   354 => x"05415f5d",
   355 => x"5b595755",
   356 => x"817b278f",
   357 => x"38767d0c",
   358 => x"77841e0c",
   359 => x"7cb00c90",
   360 => x"3d0d0480",
   361 => x"c7a80855",
   362 => x"ffba39ff",
   363 => x"3d0d80c7",
   364 => x"b0335170",
   365 => x"a73880c0",
   366 => x"80087008",
   367 => x"52527080",
   368 => x"2e943884",
   369 => x"1280c080",
   370 => x"0c702d80",
   371 => x"c0800870",
   372 => x"08525270",
   373 => x"ee38810b",
   374 => x"80c7b034",
   375 => x"833d0d04",
   376 => x"04803d0d",
   377 => x"0b0b80c7",
   378 => x"a008802e",
   379 => x"8e380b0b",
   380 => x"0b0b800b",
   381 => x"802e0981",
   382 => x"06853882",
   383 => x"3d0d040b",
   384 => x"0b80c7a0",
   385 => x"510b0b0b",
   386 => x"f3f63f82",
   387 => x"3d0d0404",
   388 => x"c008b00c",
   389 => x"04803d0d",
   390 => x"80c10b81",
   391 => x"97943480",
   392 => x"0b8199ac",
   393 => x"0c70b00c",
   394 => x"823d0d04",
   395 => x"ff3d0d80",
   396 => x"0b819794",
   397 => x"33525270",
   398 => x"80c12e99",
   399 => x"38718199",
   400 => x"ac080781",
   401 => x"99ac0c80",
   402 => x"c20b8197",
   403 => x"983470b0",
   404 => x"0c833d0d",
   405 => x"04810b81",
   406 => x"99ac0807",
   407 => x"8199ac0c",
   408 => x"80c20b81",
   409 => x"97983470",
   410 => x"b00c833d",
   411 => x"0d04fd3d",
   412 => x"0d757008",
   413 => x"8a055353",
   414 => x"81979433",
   415 => x"517080c1",
   416 => x"2e8b3873",
   417 => x"f33870b0",
   418 => x"0c853d0d",
   419 => x"04ff1270",
   420 => x"81979008",
   421 => x"31740cb0",
   422 => x"0c853d0d",
   423 => x"04fc3d0d",
   424 => x"8197bc08",
   425 => x"5574802e",
   426 => x"8c387675",
   427 => x"08710c81",
   428 => x"97bc0856",
   429 => x"548c1553",
   430 => x"81979008",
   431 => x"528a518c",
   432 => x"a33f73b0",
   433 => x"0c863d0d",
   434 => x"04fb3d0d",
   435 => x"77700856",
   436 => x"56b05381",
   437 => x"97bc0852",
   438 => x"745198c0",
   439 => x"3f850b8c",
   440 => x"170c850b",
   441 => x"8c160c75",
   442 => x"08750c81",
   443 => x"97bc0854",
   444 => x"73802e8a",
   445 => x"38730875",
   446 => x"0c8197bc",
   447 => x"08548c14",
   448 => x"53819790",
   449 => x"08528a51",
   450 => x"8bda3f84",
   451 => x"1508ad38",
   452 => x"860b8c16",
   453 => x"0c881552",
   454 => x"88160851",
   455 => x"8ae63f81",
   456 => x"97bc0870",
   457 => x"08760c54",
   458 => x"8c157054",
   459 => x"548a5273",
   460 => x"08518bb0",
   461 => x"3f73b00c",
   462 => x"873d0d04",
   463 => x"750854b0",
   464 => x"53735275",
   465 => x"5197d53f",
   466 => x"73b00c87",
   467 => x"3d0d04f3",
   468 => x"3d0d88bd",
   469 => x"0bff880c",
   470 => x"8196a80b",
   471 => x"8196dc0c",
   472 => x"8196e00b",
   473 => x"8197bc0c",
   474 => x"8196a80b",
   475 => x"8196e00c",
   476 => x"800b8196",
   477 => x"e00b8405",
   478 => x"0c820b81",
   479 => x"96e00b88",
   480 => x"050ca80b",
   481 => x"8196e00b",
   482 => x"8c050c9f",
   483 => x"53b3e052",
   484 => x"8196f051",
   485 => x"97863f9f",
   486 => x"53b48052",
   487 => x"81998c51",
   488 => x"96fa3f8a",
   489 => x"0b80d4f4",
   490 => x"0cbea451",
   491 => x"8da63fb4",
   492 => x"a0518da0",
   493 => x"3fbea451",
   494 => x"8d9a3f80",
   495 => x"c0880880",
   496 => x"2e87d238",
   497 => x"b4d0518d",
   498 => x"8b3fbea4",
   499 => x"518d853f",
   500 => x"80c08408",
   501 => x"52b4fc51",
   502 => x"8cfa3fc0",
   503 => x"0880c894",
   504 => x"0c815880",
   505 => x"0b80c084",
   506 => x"082582d0",
   507 => x"388c3d5b",
   508 => x"80c10b81",
   509 => x"97943481",
   510 => x"0b8199ac",
   511 => x"0c80c20b",
   512 => x"81979834",
   513 => x"825c835a",
   514 => x"9f53b5ac",
   515 => x"5281979c",
   516 => x"5196893f",
   517 => x"815d800b",
   518 => x"81979c53",
   519 => x"81998c52",
   520 => x"558ae53f",
   521 => x"b008752e",
   522 => x"09810683",
   523 => x"38815574",
   524 => x"8199ac0c",
   525 => x"7b705755",
   526 => x"748325a0",
   527 => x"38741010",
   528 => x"15fd055e",
   529 => x"8f3dfc05",
   530 => x"53835275",
   531 => x"5189953f",
   532 => x"811c705d",
   533 => x"70575583",
   534 => x"7524e238",
   535 => x"7d547453",
   536 => x"80c89852",
   537 => x"8197c451",
   538 => x"898a3f81",
   539 => x"97bc0870",
   540 => x"085757b0",
   541 => x"53765275",
   542 => x"5195a13f",
   543 => x"850b8c18",
   544 => x"0c850b8c",
   545 => x"170c7608",
   546 => x"760c8197",
   547 => x"bc085574",
   548 => x"802e8a38",
   549 => x"7408760c",
   550 => x"8197bc08",
   551 => x"558c1553",
   552 => x"81979008",
   553 => x"528a5188",
   554 => x"bb3f8416",
   555 => x"08878e38",
   556 => x"860b8c17",
   557 => x"0c881652",
   558 => x"88170851",
   559 => x"87c63f81",
   560 => x"97bc0870",
   561 => x"08770c55",
   562 => x"8c167054",
   563 => x"578a5276",
   564 => x"08518890",
   565 => x"3f80c10b",
   566 => x"81979833",
   567 => x"56567575",
   568 => x"26a23880",
   569 => x"c3527551",
   570 => x"88f43fb0",
   571 => x"087d2e86",
   572 => x"9f388116",
   573 => x"7081ff06",
   574 => x"81979833",
   575 => x"57575774",
   576 => x"7627e038",
   577 => x"797c297e",
   578 => x"70723570",
   579 => x"5f727231",
   580 => x"70872972",
   581 => x"3153538a",
   582 => x"05819794",
   583 => x"33819790",
   584 => x"085a5a52",
   585 => x"5b557680",
   586 => x"c12e86a9",
   587 => x"3878f738",
   588 => x"81185880",
   589 => x"c0840878",
   590 => x"25fdb538",
   591 => x"c0088196",
   592 => x"d80cb5cc",
   593 => x"518a8d3f",
   594 => x"bea4518a",
   595 => x"873fb5dc",
   596 => x"518a813f",
   597 => x"bea45189",
   598 => x"fb3f8197",
   599 => x"900852b6",
   600 => x"945189f0",
   601 => x"3f8552b6",
   602 => x"b05189e8",
   603 => x"3f8199ac",
   604 => x"0852b6cc",
   605 => x"5189dd3f",
   606 => x"8152b6b0",
   607 => x"5189d53f",
   608 => x"81979433",
   609 => x"52b6e851",
   610 => x"89ca3f80",
   611 => x"c152b784",
   612 => x"5189c13f",
   613 => x"81979833",
   614 => x"52b7a051",
   615 => x"89b63f80",
   616 => x"c252b784",
   617 => x"5189ad3f",
   618 => x"8197e408",
   619 => x"52b7bc51",
   620 => x"89a23f87",
   621 => x"52b6b051",
   622 => x"899a3f80",
   623 => x"d4f40852",
   624 => x"b7d85189",
   625 => x"8f3fb7f4",
   626 => x"5189893f",
   627 => x"b8a05189",
   628 => x"833f8197",
   629 => x"bc087008",
   630 => x"5357b8ac",
   631 => x"5188f53f",
   632 => x"b8c85188",
   633 => x"ef3f8197",
   634 => x"bc088411",
   635 => x"08535bb8",
   636 => x"fc5188e0",
   637 => x"3f8052b6",
   638 => x"b05188d8",
   639 => x"3f8197bc",
   640 => x"08881108",
   641 => x"5358b998",
   642 => x"5188c93f",
   643 => x"8252b6b0",
   644 => x"5188c13f",
   645 => x"8197bc08",
   646 => x"8c110853",
   647 => x"59b9b451",
   648 => x"88b23f91",
   649 => x"52b6b051",
   650 => x"88aa3f81",
   651 => x"97bc0890",
   652 => x"0552b9d0",
   653 => x"51889d3f",
   654 => x"b9ec5188",
   655 => x"973fbaa4",
   656 => x"5188913f",
   657 => x"8196dc08",
   658 => x"70085355",
   659 => x"b8ac5188",
   660 => x"833fbab8",
   661 => x"5187fd3f",
   662 => x"8196dc08",
   663 => x"84110853",
   664 => x"56b8fc51",
   665 => x"87ee3f80",
   666 => x"52b6b051",
   667 => x"87e63f81",
   668 => x"96dc0888",
   669 => x"11085357",
   670 => x"b9985187",
   671 => x"d73f8152",
   672 => x"b6b05187",
   673 => x"cf3f8196",
   674 => x"dc088c11",
   675 => x"08535bb9",
   676 => x"b45187c0",
   677 => x"3f9252b6",
   678 => x"b05187b8",
   679 => x"3f8196dc",
   680 => x"08900552",
   681 => x"b9d05187",
   682 => x"ab3fb9ec",
   683 => x"5187a53f",
   684 => x"7b52baf8",
   685 => x"51879d3f",
   686 => x"8552b6b0",
   687 => x"5187953f",
   688 => x"7952bb94",
   689 => x"51878d3f",
   690 => x"8d52b6b0",
   691 => x"5187853f",
   692 => x"7d52bbb0",
   693 => x"5186fd3f",
   694 => x"8752b6b0",
   695 => x"5186f53f",
   696 => x"7c52bbcc",
   697 => x"5186ed3f",
   698 => x"8152b6b0",
   699 => x"5186e53f",
   700 => x"81998c52",
   701 => x"bbe85186",
   702 => x"db3fbc84",
   703 => x"5186d53f",
   704 => x"81979c52",
   705 => x"bcbc5186",
   706 => x"cb3fbcd8",
   707 => x"5186c53f",
   708 => x"bea45186",
   709 => x"bf3f8196",
   710 => x"d80880c8",
   711 => x"94083170",
   712 => x"80c8900c",
   713 => x"52bd9051",
   714 => x"86aa3f80",
   715 => x"c8900856",
   716 => x"80f77625",
   717 => x"80e53880",
   718 => x"c0840870",
   719 => x"7787e829",
   720 => x"3580c888",
   721 => x"0c767187",
   722 => x"e8293580",
   723 => x"c88c0c76",
   724 => x"7184b929",
   725 => x"358197c0",
   726 => x"0c5abda0",
   727 => x"5185f53f",
   728 => x"80c88808",
   729 => x"52bdd051",
   730 => x"85ea3fbd",
   731 => x"d85185e4",
   732 => x"3f80c88c",
   733 => x"0852bdd0",
   734 => x"5185d93f",
   735 => x"8197c008",
   736 => x"52be8851",
   737 => x"85ce3fbe",
   738 => x"a45185c8",
   739 => x"3f800bb0",
   740 => x"0c8f3d0d",
   741 => x"04bea851",
   742 => x"f8ad39be",
   743 => x"d85185b4",
   744 => x"3fbf9051",
   745 => x"85ae3fbe",
   746 => x"a45185a8",
   747 => x"3f80c890",
   748 => x"0880c084",
   749 => x"08707287",
   750 => x"e8293580",
   751 => x"c8880c71",
   752 => x"7187e829",
   753 => x"3580c88c",
   754 => x"0c717184",
   755 => x"b9293581",
   756 => x"97c00c5b",
   757 => x"56bda051",
   758 => x"84fa3f80",
   759 => x"c8880852",
   760 => x"bdd05184",
   761 => x"ef3fbdd8",
   762 => x"5184e93f",
   763 => x"80c88c08",
   764 => x"52bdd051",
   765 => x"84de3f81",
   766 => x"97c00852",
   767 => x"be885184",
   768 => x"d33fbea4",
   769 => x"5184cd3f",
   770 => x"800bb00c",
   771 => x"8f3d0d04",
   772 => x"8f3df805",
   773 => x"52805180",
   774 => x"eb3f9f53",
   775 => x"bfb05281",
   776 => x"979c518d",
   777 => x"f73f7778",
   778 => x"8197900c",
   779 => x"81177081",
   780 => x"ff068197",
   781 => x"98335858",
   782 => x"585af9c3",
   783 => x"39760856",
   784 => x"b0537552",
   785 => x"76518dd4",
   786 => x"3f80c10b",
   787 => x"81979833",
   788 => x"5656f98a",
   789 => x"39ff1570",
   790 => x"77317c0c",
   791 => x"59800b81",
   792 => x"19595980",
   793 => x"c0840878",
   794 => x"25f78538",
   795 => x"f9ce39ff",
   796 => x"3d0d7382",
   797 => x"32703070",
   798 => x"72078025",
   799 => x"b00c5252",
   800 => x"833d0d04",
   801 => x"fe3d0d74",
   802 => x"76715354",
   803 => x"5271822e",
   804 => x"83388351",
   805 => x"71812e9a",
   806 => x"38817226",
   807 => x"9f387182",
   808 => x"2eb83871",
   809 => x"842ea938",
   810 => x"70730c70",
   811 => x"b00c843d",
   812 => x"0d0480e4",
   813 => x"0b819790",
   814 => x"08258b38",
   815 => x"80730c70",
   816 => x"b00c843d",
   817 => x"0d048373",
   818 => x"0c70b00c",
   819 => x"843d0d04",
   820 => x"82730c70",
   821 => x"b00c843d",
   822 => x"0d048173",
   823 => x"0c70b00c",
   824 => x"843d0d04",
   825 => x"803d0d74",
   826 => x"74148205",
   827 => x"710cb00c",
   828 => x"823d0d04",
   829 => x"f73d0d7b",
   830 => x"7d7f6185",
   831 => x"1270822b",
   832 => x"75117074",
   833 => x"71708405",
   834 => x"530c5a5a",
   835 => x"5d5b760c",
   836 => x"7980f818",
   837 => x"0c798612",
   838 => x"5257585a",
   839 => x"5a767624",
   840 => x"993876b3",
   841 => x"29822b79",
   842 => x"11515376",
   843 => x"73708405",
   844 => x"550c8114",
   845 => x"54757425",
   846 => x"f2387681",
   847 => x"cc2919fc",
   848 => x"11088105",
   849 => x"fc120c7a",
   850 => x"1970089f",
   851 => x"a0130c58",
   852 => x"56850b81",
   853 => x"97900c75",
   854 => x"b00c8b3d",
   855 => x"0d04fe3d",
   856 => x"0d029305",
   857 => x"33518002",
   858 => x"84059705",
   859 => x"33545270",
   860 => x"732e8838",
   861 => x"71b00c84",
   862 => x"3d0d0470",
   863 => x"81979434",
   864 => x"810bb00c",
   865 => x"843d0d04",
   866 => x"f83d0d7a",
   867 => x"7c595682",
   868 => x"0b831955",
   869 => x"55741670",
   870 => x"3375335b",
   871 => x"51537279",
   872 => x"2e80c638",
   873 => x"80c10b81",
   874 => x"16811656",
   875 => x"56578275",
   876 => x"25e338ff",
   877 => x"a9177081",
   878 => x"ff065559",
   879 => x"73822683",
   880 => x"38875581",
   881 => x"537680d2",
   882 => x"2e983877",
   883 => x"5275518b",
   884 => x"e43f8053",
   885 => x"72b00825",
   886 => x"89388715",
   887 => x"8197900c",
   888 => x"815372b0",
   889 => x"0c8a3d0d",
   890 => x"04728197",
   891 => x"94348275",
   892 => x"25ffa238",
   893 => x"ffbd39fe",
   894 => x"3d0d7470",
   895 => x"337081ff",
   896 => x"06535353",
   897 => x"70802ea7",
   898 => x"38ff8408",
   899 => x"70882a70",
   900 => x"81065151",
   901 => x"5170802e",
   902 => x"f0387181",
   903 => x"ff068114",
   904 => x"54ff840c",
   905 => x"72337081",
   906 => x"ff065252",
   907 => x"70db3884",
   908 => x"3d0d04ff",
   909 => x"3d0d028f",
   910 => x"053352ff",
   911 => x"84087088",
   912 => x"2a708106",
   913 => x"51515170",
   914 => x"802ef038",
   915 => x"71ff840c",
   916 => x"833d0d04",
   917 => x"f53d0d8e",
   918 => x"3d707084",
   919 => x"0552089c",
   920 => x"b35b555b",
   921 => x"80747081",
   922 => x"05563375",
   923 => x"5a545772",
   924 => x"772ebe38",
   925 => x"72a52e09",
   926 => x"810680c5",
   927 => x"38777081",
   928 => x"05593353",
   929 => x"7280e42e",
   930 => x"81b63872",
   931 => x"80e42480",
   932 => x"c6387280",
   933 => x"e32ea138",
   934 => x"8052a551",
   935 => x"782d8052",
   936 => x"7251782d",
   937 => x"82175777",
   938 => x"70810559",
   939 => x"335372c4",
   940 => x"3876b00c",
   941 => x"8d3d0d04",
   942 => x"7a841c83",
   943 => x"1233555c",
   944 => x"56805272",
   945 => x"51782d81",
   946 => x"17787081",
   947 => x"055a3354",
   948 => x"5772ffa0",
   949 => x"38db3972",
   950 => x"80f32e09",
   951 => x"8106ffb8",
   952 => x"387a841c",
   953 => x"7108585c",
   954 => x"54807633",
   955 => x"5b557975",
   956 => x"2e8d3881",
   957 => x"15701770",
   958 => x"33555b55",
   959 => x"72f538ff",
   960 => x"15548075",
   961 => x"25ffa038",
   962 => x"75708105",
   963 => x"57335380",
   964 => x"52725178",
   965 => x"2d811774",
   966 => x"ff165656",
   967 => x"57807525",
   968 => x"ff853875",
   969 => x"70810557",
   970 => x"33538052",
   971 => x"7251782d",
   972 => x"811774ff",
   973 => x"16565657",
   974 => x"748024cc",
   975 => x"38fee839",
   976 => x"7a841c71",
   977 => x"088199c0",
   978 => x"0b80c7b4",
   979 => x"545d565c",
   980 => x"55805673",
   981 => x"762e0981",
   982 => x"06b838b0",
   983 => x"0b80c7b4",
   984 => x"34811555",
   985 => x"ff155574",
   986 => x"337a7081",
   987 => x"055c3481",
   988 => x"16567480",
   989 => x"c7b42e09",
   990 => x"8106e938",
   991 => x"807a3475",
   992 => x"8199c00b",
   993 => x"ff125657",
   994 => x"55748024",
   995 => x"fefa38fe",
   996 => x"9639738f",
   997 => x"06bfd005",
   998 => x"53723375",
   999 => x"70810557",
  1000 => x"3473842a",
  1001 => x"5473eb38",
  1002 => x"7480c7b4",
  1003 => x"2ece38ff",
  1004 => x"15557433",
  1005 => x"7a708105",
  1006 => x"5c348116",
  1007 => x"567480c7",
  1008 => x"b42effb8",
  1009 => x"38ff9d39",
  1010 => x"bc0802bc",
  1011 => x"0cf53d0d",
  1012 => x"bc089405",
  1013 => x"089d38bc",
  1014 => x"088c0508",
  1015 => x"bc089005",
  1016 => x"08bc0888",
  1017 => x"05085856",
  1018 => x"5473760c",
  1019 => x"7484170c",
  1020 => x"81bf3980",
  1021 => x"0bbc08f0",
  1022 => x"050c800b",
  1023 => x"bc08f405",
  1024 => x"0cbc088c",
  1025 => x"0508bc08",
  1026 => x"90050856",
  1027 => x"5473bc08",
  1028 => x"f0050c74",
  1029 => x"bc08f405",
  1030 => x"0cbc08f8",
  1031 => x"05bc08f0",
  1032 => x"05565688",
  1033 => x"70547553",
  1034 => x"76525485",
  1035 => x"ef3fa00b",
  1036 => x"bc089405",
  1037 => x"0831bc08",
  1038 => x"ec050cbc",
  1039 => x"08ec0508",
  1040 => x"80249d38",
  1041 => x"800bbc08",
  1042 => x"f4050cbc",
  1043 => x"08ec0508",
  1044 => x"30bc08fc",
  1045 => x"0508712b",
  1046 => x"bc08f005",
  1047 => x"0c54b939",
  1048 => x"bc08fc05",
  1049 => x"08bc08ec",
  1050 => x"05082abc",
  1051 => x"08e8050c",
  1052 => x"bc08fc05",
  1053 => x"08bc0894",
  1054 => x"05082bbc",
  1055 => x"08f4050c",
  1056 => x"bc08f805",
  1057 => x"08bc0894",
  1058 => x"05082b70",
  1059 => x"bc08e805",
  1060 => x"0807bc08",
  1061 => x"f0050c54",
  1062 => x"bc08f005",
  1063 => x"08bc08f4",
  1064 => x"0508bc08",
  1065 => x"88050858",
  1066 => x"56547376",
  1067 => x"0c748417",
  1068 => x"0cbc0888",
  1069 => x"0508b00c",
  1070 => x"8d3d0dbc",
  1071 => x"0c04bc08",
  1072 => x"02bc0cf9",
  1073 => x"3d0d800b",
  1074 => x"bc08fc05",
  1075 => x"0cbc0888",
  1076 => x"05088025",
  1077 => x"ab38bc08",
  1078 => x"88050830",
  1079 => x"bc088805",
  1080 => x"0c800bbc",
  1081 => x"08f4050c",
  1082 => x"bc08fc05",
  1083 => x"08883881",
  1084 => x"0bbc08f4",
  1085 => x"050cbc08",
  1086 => x"f40508bc",
  1087 => x"08fc050c",
  1088 => x"bc088c05",
  1089 => x"088025ab",
  1090 => x"38bc088c",
  1091 => x"050830bc",
  1092 => x"088c050c",
  1093 => x"800bbc08",
  1094 => x"f0050cbc",
  1095 => x"08fc0508",
  1096 => x"8838810b",
  1097 => x"bc08f005",
  1098 => x"0cbc08f0",
  1099 => x"0508bc08",
  1100 => x"fc050c80",
  1101 => x"53bc088c",
  1102 => x"050852bc",
  1103 => x"08880508",
  1104 => x"5181a73f",
  1105 => x"b00870bc",
  1106 => x"08f8050c",
  1107 => x"54bc08fc",
  1108 => x"0508802e",
  1109 => x"8c38bc08",
  1110 => x"f8050830",
  1111 => x"bc08f805",
  1112 => x"0cbc08f8",
  1113 => x"050870b0",
  1114 => x"0c54893d",
  1115 => x"0dbc0c04",
  1116 => x"bc0802bc",
  1117 => x"0cfb3d0d",
  1118 => x"800bbc08",
  1119 => x"fc050cbc",
  1120 => x"08880508",
  1121 => x"80259338",
  1122 => x"bc088805",
  1123 => x"0830bc08",
  1124 => x"88050c81",
  1125 => x"0bbc08fc",
  1126 => x"050cbc08",
  1127 => x"8c050880",
  1128 => x"258c38bc",
  1129 => x"088c0508",
  1130 => x"30bc088c",
  1131 => x"050c8153",
  1132 => x"bc088c05",
  1133 => x"0852bc08",
  1134 => x"88050851",
  1135 => x"ad3fb008",
  1136 => x"70bc08f8",
  1137 => x"050c54bc",
  1138 => x"08fc0508",
  1139 => x"802e8c38",
  1140 => x"bc08f805",
  1141 => x"0830bc08",
  1142 => x"f8050cbc",
  1143 => x"08f80508",
  1144 => x"70b00c54",
  1145 => x"873d0dbc",
  1146 => x"0c04bc08",
  1147 => x"02bc0cfd",
  1148 => x"3d0d810b",
  1149 => x"bc08fc05",
  1150 => x"0c800bbc",
  1151 => x"08f8050c",
  1152 => x"bc088c05",
  1153 => x"08bc0888",
  1154 => x"050827ac",
  1155 => x"38bc08fc",
  1156 => x"0508802e",
  1157 => x"a338800b",
  1158 => x"bc088c05",
  1159 => x"08249938",
  1160 => x"bc088c05",
  1161 => x"0810bc08",
  1162 => x"8c050cbc",
  1163 => x"08fc0508",
  1164 => x"10bc08fc",
  1165 => x"050cc939",
  1166 => x"bc08fc05",
  1167 => x"08802e80",
  1168 => x"c938bc08",
  1169 => x"8c0508bc",
  1170 => x"08880508",
  1171 => x"26a138bc",
  1172 => x"08880508",
  1173 => x"bc088c05",
  1174 => x"0831bc08",
  1175 => x"88050cbc",
  1176 => x"08f80508",
  1177 => x"bc08fc05",
  1178 => x"0807bc08",
  1179 => x"f8050cbc",
  1180 => x"08fc0508",
  1181 => x"812abc08",
  1182 => x"fc050cbc",
  1183 => x"088c0508",
  1184 => x"812abc08",
  1185 => x"8c050cff",
  1186 => x"af39bc08",
  1187 => x"90050880",
  1188 => x"2e8f38bc",
  1189 => x"08880508",
  1190 => x"70bc08f4",
  1191 => x"050c518d",
  1192 => x"39bc08f8",
  1193 => x"050870bc",
  1194 => x"08f4050c",
  1195 => x"51bc08f4",
  1196 => x"0508b00c",
  1197 => x"853d0dbc",
  1198 => x"0c04bc08",
  1199 => x"02bc0cff",
  1200 => x"3d0d800b",
  1201 => x"bc08fc05",
  1202 => x"0cbc0888",
  1203 => x"05088106",
  1204 => x"ff117009",
  1205 => x"70bc088c",
  1206 => x"050806bc",
  1207 => x"08fc0508",
  1208 => x"11bc08fc",
  1209 => x"050cbc08",
  1210 => x"88050881",
  1211 => x"2abc0888",
  1212 => x"050cbc08",
  1213 => x"8c050810",
  1214 => x"bc088c05",
  1215 => x"0c515151",
  1216 => x"51bc0888",
  1217 => x"0508802e",
  1218 => x"8438ffbd",
  1219 => x"39bc08fc",
  1220 => x"050870b0",
  1221 => x"0c51833d",
  1222 => x"0dbc0c04",
  1223 => x"fc3d0d76",
  1224 => x"70797b55",
  1225 => x"5555558f",
  1226 => x"72278c38",
  1227 => x"72750783",
  1228 => x"06517080",
  1229 => x"2ea738ff",
  1230 => x"125271ff",
  1231 => x"2e983872",
  1232 => x"70810554",
  1233 => x"33747081",
  1234 => x"055634ff",
  1235 => x"125271ff",
  1236 => x"2e098106",
  1237 => x"ea3874b0",
  1238 => x"0c863d0d",
  1239 => x"04745172",
  1240 => x"70840554",
  1241 => x"08717084",
  1242 => x"05530c72",
  1243 => x"70840554",
  1244 => x"08717084",
  1245 => x"05530c72",
  1246 => x"70840554",
  1247 => x"08717084",
  1248 => x"05530c72",
  1249 => x"70840554",
  1250 => x"08717084",
  1251 => x"05530cf0",
  1252 => x"1252718f",
  1253 => x"26c93883",
  1254 => x"72279538",
  1255 => x"72708405",
  1256 => x"54087170",
  1257 => x"8405530c",
  1258 => x"fc125271",
  1259 => x"8326ed38",
  1260 => x"7054ff83",
  1261 => x"39fb3d0d",
  1262 => x"77797072",
  1263 => x"07830653",
  1264 => x"54527093",
  1265 => x"38717373",
  1266 => x"08545654",
  1267 => x"7173082e",
  1268 => x"80c43873",
  1269 => x"75545271",
  1270 => x"337081ff",
  1271 => x"06525470",
  1272 => x"802e9d38",
  1273 => x"72335570",
  1274 => x"752e0981",
  1275 => x"06953881",
  1276 => x"12811471",
  1277 => x"337081ff",
  1278 => x"06545654",
  1279 => x"5270e538",
  1280 => x"72335573",
  1281 => x"81ff0675",
  1282 => x"81ff0671",
  1283 => x"7131b00c",
  1284 => x"5252873d",
  1285 => x"0d047109",
  1286 => x"70f7fbfd",
  1287 => x"ff140670",
  1288 => x"f8848281",
  1289 => x"80065151",
  1290 => x"51709738",
  1291 => x"84148416",
  1292 => x"71085456",
  1293 => x"54717508",
  1294 => x"2edc3873",
  1295 => x"755452ff",
  1296 => x"9639800b",
  1297 => x"b00c873d",
  1298 => x"0d04fd3d",
  1299 => x"0d800bbf",
  1300 => x"f8085454",
  1301 => x"72812e9b",
  1302 => x"387380c8",
  1303 => x"840ce185",
  1304 => x"3fdf9d3f",
  1305 => x"80c08c52",
  1306 => x"8151e5e3",
  1307 => x"3fb00851",
  1308 => x"879b3f72",
  1309 => x"80c8840c",
  1310 => x"e0eb3fdf",
  1311 => x"833f80c0",
  1312 => x"8c528151",
  1313 => x"e5c93fb0",
  1314 => x"08518781",
  1315 => x"3f00ff39",
  1316 => x"00ff39f5",
  1317 => x"3d0d7e60",
  1318 => x"80c88408",
  1319 => x"705b585b",
  1320 => x"5b7580c2",
  1321 => x"38777a25",
  1322 => x"a138771b",
  1323 => x"70337081",
  1324 => x"ff065858",
  1325 => x"59758a2e",
  1326 => x"98387681",
  1327 => x"ff0651e0",
  1328 => x"833f8118",
  1329 => x"58797824",
  1330 => x"e13879b0",
  1331 => x"0c8d3d0d",
  1332 => x"048d51df",
  1333 => x"ef3f7833",
  1334 => x"7081ff06",
  1335 => x"5257dfe4",
  1336 => x"3f811858",
  1337 => x"e0397955",
  1338 => x"7a547d53",
  1339 => x"85528d3d",
  1340 => x"fc0551de",
  1341 => x"cc3fb008",
  1342 => x"56868b3f",
  1343 => x"7bb0080c",
  1344 => x"75b00c8d",
  1345 => x"3d0d04f6",
  1346 => x"3d0d7d7f",
  1347 => x"80c88408",
  1348 => x"705b585a",
  1349 => x"5a7580c1",
  1350 => x"38777925",
  1351 => x"b338deff",
  1352 => x"3fb00881",
  1353 => x"ff06708d",
  1354 => x"32703070",
  1355 => x"9f2a5151",
  1356 => x"5757768a",
  1357 => x"2e80c338",
  1358 => x"75802ebe",
  1359 => x"38771a56",
  1360 => x"76763476",
  1361 => x"51defd3f",
  1362 => x"81185878",
  1363 => x"7824cf38",
  1364 => x"775675b0",
  1365 => x"0c8c3d0d",
  1366 => x"04785579",
  1367 => x"547c5384",
  1368 => x"528c3dfc",
  1369 => x"0551ddd9",
  1370 => x"3fb00856",
  1371 => x"85983f7a",
  1372 => x"b0080c75",
  1373 => x"b00c8c3d",
  1374 => x"0d04771a",
  1375 => x"568a7634",
  1376 => x"8118588d",
  1377 => x"51debd3f",
  1378 => x"8a51deb8",
  1379 => x"3f7756c2",
  1380 => x"39f93d0d",
  1381 => x"795780c8",
  1382 => x"8408802e",
  1383 => x"ac387651",
  1384 => x"879e3f7b",
  1385 => x"567a55b0",
  1386 => x"08810554",
  1387 => x"76538252",
  1388 => x"893dfc05",
  1389 => x"51dd8a3f",
  1390 => x"b0085784",
  1391 => x"c93f77b0",
  1392 => x"080c76b0",
  1393 => x"0c893d0d",
  1394 => x"0484bb3f",
  1395 => x"850bb008",
  1396 => x"0cff0bb0",
  1397 => x"0c893d0d",
  1398 => x"04fb3d0d",
  1399 => x"80c88408",
  1400 => x"70565473",
  1401 => x"883874b0",
  1402 => x"0c873d0d",
  1403 => x"04775383",
  1404 => x"52873dfc",
  1405 => x"0551dcc9",
  1406 => x"3fb00854",
  1407 => x"84883f75",
  1408 => x"b0080c73",
  1409 => x"b00c873d",
  1410 => x"0d04ff0b",
  1411 => x"b00c04fb",
  1412 => x"3d0d7755",
  1413 => x"80c88408",
  1414 => x"802ea838",
  1415 => x"745186a0",
  1416 => x"3fb00881",
  1417 => x"05547453",
  1418 => x"8752873d",
  1419 => x"fc0551dc",
  1420 => x"903fb008",
  1421 => x"5583cf3f",
  1422 => x"75b0080c",
  1423 => x"74b00c87",
  1424 => x"3d0d0483",
  1425 => x"c13f850b",
  1426 => x"b0080cff",
  1427 => x"0bb00c87",
  1428 => x"3d0d04fa",
  1429 => x"3d0d80c8",
  1430 => x"8408802e",
  1431 => x"a2387a55",
  1432 => x"79547853",
  1433 => x"8652883d",
  1434 => x"fc0551db",
  1435 => x"d43fb008",
  1436 => x"5683933f",
  1437 => x"76b0080c",
  1438 => x"75b00c88",
  1439 => x"3d0d0483",
  1440 => x"853f9d0b",
  1441 => x"b0080cff",
  1442 => x"0bb00c88",
  1443 => x"3d0d04fb",
  1444 => x"3d0d7779",
  1445 => x"56568070",
  1446 => x"54547375",
  1447 => x"259f3874",
  1448 => x"101010f8",
  1449 => x"05527216",
  1450 => x"70337074",
  1451 => x"2b760781",
  1452 => x"16f81656",
  1453 => x"56565151",
  1454 => x"747324ea",
  1455 => x"3873b00c",
  1456 => x"873d0d04",
  1457 => x"fc3d0d76",
  1458 => x"785555bc",
  1459 => x"53805273",
  1460 => x"5183de3f",
  1461 => x"84527451",
  1462 => x"ffb53fb0",
  1463 => x"08742384",
  1464 => x"52841551",
  1465 => x"ffa93fb0",
  1466 => x"08821523",
  1467 => x"84528815",
  1468 => x"51ff9c3f",
  1469 => x"b0088415",
  1470 => x"0c84528c",
  1471 => x"1551ff8f",
  1472 => x"3fb00888",
  1473 => x"15238452",
  1474 => x"901551ff",
  1475 => x"823fb008",
  1476 => x"8a152384",
  1477 => x"52941551",
  1478 => x"fef53fb0",
  1479 => x"088c1523",
  1480 => x"84529815",
  1481 => x"51fee83f",
  1482 => x"b0088e15",
  1483 => x"2388529c",
  1484 => x"1551fedb",
  1485 => x"3fb00890",
  1486 => x"150c863d",
  1487 => x"0d04e93d",
  1488 => x"0d6a80c8",
  1489 => x"84085757",
  1490 => x"75933880",
  1491 => x"c0800b84",
  1492 => x"180c75ac",
  1493 => x"180c75b0",
  1494 => x"0c993d0d",
  1495 => x"04893d70",
  1496 => x"556a5455",
  1497 => x"8a52993d",
  1498 => x"ffbc0551",
  1499 => x"d9d33fb0",
  1500 => x"08775375",
  1501 => x"5256fecc",
  1502 => x"3f818b3f",
  1503 => x"77b0080c",
  1504 => x"75b00c99",
  1505 => x"3d0d04e9",
  1506 => x"3d0d6957",
  1507 => x"80c88408",
  1508 => x"802eb538",
  1509 => x"765183a8",
  1510 => x"3f893d70",
  1511 => x"56b00881",
  1512 => x"05557754",
  1513 => x"568f5299",
  1514 => x"3dffbc05",
  1515 => x"51d9923f",
  1516 => x"b0086b53",
  1517 => x"765257fe",
  1518 => x"8b3f80ca",
  1519 => x"3f77b008",
  1520 => x"0c76b00c",
  1521 => x"993d0d04",
  1522 => x"bd3f850b",
  1523 => x"b0080cff",
  1524 => x"0bb00c99",
  1525 => x"3d0d04fc",
  1526 => x"3d0d8154",
  1527 => x"80c88408",
  1528 => x"883873b0",
  1529 => x"0c863d0d",
  1530 => x"04765397",
  1531 => x"b952863d",
  1532 => x"fc0551d8",
  1533 => x"cc3fb008",
  1534 => x"548c3f74",
  1535 => x"b0080c73",
  1536 => x"b00c863d",
  1537 => x"0d0480c0",
  1538 => x"9008b00c",
  1539 => x"04f73d0d",
  1540 => x"7b80c090",
  1541 => x"0882c811",
  1542 => x"085a545a",
  1543 => x"77802e80",
  1544 => x"da388188",
  1545 => x"18841908",
  1546 => x"ff058171",
  1547 => x"2b595559",
  1548 => x"80742480",
  1549 => x"ea388074",
  1550 => x"24b53873",
  1551 => x"822b7811",
  1552 => x"88055656",
  1553 => x"81801908",
  1554 => x"77065372",
  1555 => x"802eb638",
  1556 => x"78167008",
  1557 => x"53537951",
  1558 => x"74085372",
  1559 => x"2dff14fc",
  1560 => x"17fc1779",
  1561 => x"812c5a57",
  1562 => x"57547380",
  1563 => x"25d63877",
  1564 => x"085877ff",
  1565 => x"ad3880c0",
  1566 => x"900853bc",
  1567 => x"1308a538",
  1568 => x"7951f889",
  1569 => x"3f740853",
  1570 => x"722dff14",
  1571 => x"fc17fc17",
  1572 => x"79812c5a",
  1573 => x"57575473",
  1574 => x"8025ffa8",
  1575 => x"38d13980",
  1576 => x"57ff9339",
  1577 => x"7251bc13",
  1578 => x"0853722d",
  1579 => x"7951f7dd",
  1580 => x"3ffc3d0d",
  1581 => x"76797102",
  1582 => x"8c059f05",
  1583 => x"33575553",
  1584 => x"55837227",
  1585 => x"8a387483",
  1586 => x"06517080",
  1587 => x"2ea238ff",
  1588 => x"125271ff",
  1589 => x"2e933873",
  1590 => x"73708105",
  1591 => x"5534ff12",
  1592 => x"5271ff2e",
  1593 => x"098106ef",
  1594 => x"3874b00c",
  1595 => x"863d0d04",
  1596 => x"7474882b",
  1597 => x"75077071",
  1598 => x"902b0751",
  1599 => x"54518f72",
  1600 => x"27a53872",
  1601 => x"71708405",
  1602 => x"530c7271",
  1603 => x"70840553",
  1604 => x"0c727170",
  1605 => x"8405530c",
  1606 => x"72717084",
  1607 => x"05530cf0",
  1608 => x"1252718f",
  1609 => x"26dd3883",
  1610 => x"72279038",
  1611 => x"72717084",
  1612 => x"05530cfc",
  1613 => x"12527183",
  1614 => x"26f23870",
  1615 => x"53ff9039",
  1616 => x"fd3d0d75",
  1617 => x"70718306",
  1618 => x"53555270",
  1619 => x"b8387170",
  1620 => x"087009f7",
  1621 => x"fbfdff12",
  1622 => x"0670f884",
  1623 => x"82818006",
  1624 => x"51515253",
  1625 => x"709d3884",
  1626 => x"13700870",
  1627 => x"09f7fbfd",
  1628 => x"ff120670",
  1629 => x"f8848281",
  1630 => x"80065151",
  1631 => x"52537080",
  1632 => x"2ee53872",
  1633 => x"52713351",
  1634 => x"70802e8a",
  1635 => x"38811270",
  1636 => x"33525270",
  1637 => x"f8387174",
  1638 => x"31b00c85",
  1639 => x"3d0d04ff",
  1640 => x"3d0d80c7",
  1641 => x"940bfc05",
  1642 => x"70085252",
  1643 => x"70ff2e91",
  1644 => x"38702dfc",
  1645 => x"12700852",
  1646 => x"5270ff2e",
  1647 => x"098106f1",
  1648 => x"38833d0d",
  1649 => x"0404d7e3",
  1650 => x"3f040000",
  1651 => x"00ffffff",
  1652 => x"ff00ffff",
  1653 => x"ffff00ff",
  1654 => x"ffffff00",
  1655 => x"00000040",
  1656 => x"44485259",
  1657 => x"53544f4e",
  1658 => x"45205052",
  1659 => x"4f475241",
  1660 => x"4d2c2053",
  1661 => x"4f4d4520",
  1662 => x"53545249",
  1663 => x"4e470000",
  1664 => x"44485259",
  1665 => x"53544f4e",
  1666 => x"45205052",
  1667 => x"4f475241",
  1668 => x"4d2c2031",
  1669 => x"27535420",
  1670 => x"53545249",
  1671 => x"4e470000",
  1672 => x"44687279",
  1673 => x"73746f6e",
  1674 => x"65204265",
  1675 => x"6e63686d",
  1676 => x"61726b2c",
  1677 => x"20566572",
  1678 => x"73696f6e",
  1679 => x"20322e31",
  1680 => x"20284c61",
  1681 => x"6e677561",
  1682 => x"67653a20",
  1683 => x"43290a00",
  1684 => x"50726f67",
  1685 => x"72616d20",
  1686 => x"636f6d70",
  1687 => x"696c6564",
  1688 => x"20776974",
  1689 => x"68202772",
  1690 => x"65676973",
  1691 => x"74657227",
  1692 => x"20617474",
  1693 => x"72696275",
  1694 => x"74650a00",
  1695 => x"45786563",
  1696 => x"7574696f",
  1697 => x"6e207374",
  1698 => x"61727473",
  1699 => x"2c202564",
  1700 => x"2072756e",
  1701 => x"73207468",
  1702 => x"726f7567",
  1703 => x"68204468",
  1704 => x"72797374",
  1705 => x"6f6e650a",
  1706 => x"00000000",
  1707 => x"44485259",
  1708 => x"53544f4e",
  1709 => x"45205052",
  1710 => x"4f475241",
  1711 => x"4d2c2032",
  1712 => x"274e4420",
  1713 => x"53545249",
  1714 => x"4e470000",
  1715 => x"45786563",
  1716 => x"7574696f",
  1717 => x"6e20656e",
  1718 => x"64730a00",
  1719 => x"46696e61",
  1720 => x"6c207661",
  1721 => x"6c756573",
  1722 => x"206f6620",
  1723 => x"74686520",
  1724 => x"76617269",
  1725 => x"61626c65",
  1726 => x"73207573",
  1727 => x"65642069",
  1728 => x"6e207468",
  1729 => x"65206265",
  1730 => x"6e63686d",
  1731 => x"61726b3a",
  1732 => x"0a000000",
  1733 => x"496e745f",
  1734 => x"476c6f62",
  1735 => x"3a202020",
  1736 => x"20202020",
  1737 => x"20202020",
  1738 => x"2025640a",
  1739 => x"00000000",
  1740 => x"20202020",
  1741 => x"20202020",
  1742 => x"73686f75",
  1743 => x"6c642062",
  1744 => x"653a2020",
  1745 => x"2025640a",
  1746 => x"00000000",
  1747 => x"426f6f6c",
  1748 => x"5f476c6f",
  1749 => x"623a2020",
  1750 => x"20202020",
  1751 => x"20202020",
  1752 => x"2025640a",
  1753 => x"00000000",
  1754 => x"43685f31",
  1755 => x"5f476c6f",
  1756 => x"623a2020",
  1757 => x"20202020",
  1758 => x"20202020",
  1759 => x"2025630a",
  1760 => x"00000000",
  1761 => x"20202020",
  1762 => x"20202020",
  1763 => x"73686f75",
  1764 => x"6c642062",
  1765 => x"653a2020",
  1766 => x"2025630a",
  1767 => x"00000000",
  1768 => x"43685f32",
  1769 => x"5f476c6f",
  1770 => x"623a2020",
  1771 => x"20202020",
  1772 => x"20202020",
  1773 => x"2025630a",
  1774 => x"00000000",
  1775 => x"4172725f",
  1776 => x"315f476c",
  1777 => x"6f625b38",
  1778 => x"5d3a2020",
  1779 => x"20202020",
  1780 => x"2025640a",
  1781 => x"00000000",
  1782 => x"4172725f",
  1783 => x"325f476c",
  1784 => x"6f625b38",
  1785 => x"5d5b375d",
  1786 => x"3a202020",
  1787 => x"2025640a",
  1788 => x"00000000",
  1789 => x"20202020",
  1790 => x"20202020",
  1791 => x"73686f75",
  1792 => x"6c642062",
  1793 => x"653a2020",
  1794 => x"204e756d",
  1795 => x"6265725f",
  1796 => x"4f665f52",
  1797 => x"756e7320",
  1798 => x"2b203130",
  1799 => x"0a000000",
  1800 => x"5074725f",
  1801 => x"476c6f62",
  1802 => x"2d3e0a00",
  1803 => x"20205074",
  1804 => x"725f436f",
  1805 => x"6d703a20",
  1806 => x"20202020",
  1807 => x"20202020",
  1808 => x"2025640a",
  1809 => x"00000000",
  1810 => x"20202020",
  1811 => x"20202020",
  1812 => x"73686f75",
  1813 => x"6c642062",
  1814 => x"653a2020",
  1815 => x"2028696d",
  1816 => x"706c656d",
  1817 => x"656e7461",
  1818 => x"74696f6e",
  1819 => x"2d646570",
  1820 => x"656e6465",
  1821 => x"6e74290a",
  1822 => x"00000000",
  1823 => x"20204469",
  1824 => x"7363723a",
  1825 => x"20202020",
  1826 => x"20202020",
  1827 => x"20202020",
  1828 => x"2025640a",
  1829 => x"00000000",
  1830 => x"2020456e",
  1831 => x"756d5f43",
  1832 => x"6f6d703a",
  1833 => x"20202020",
  1834 => x"20202020",
  1835 => x"2025640a",
  1836 => x"00000000",
  1837 => x"2020496e",
  1838 => x"745f436f",
  1839 => x"6d703a20",
  1840 => x"20202020",
  1841 => x"20202020",
  1842 => x"2025640a",
  1843 => x"00000000",
  1844 => x"20205374",
  1845 => x"725f436f",
  1846 => x"6d703a20",
  1847 => x"20202020",
  1848 => x"20202020",
  1849 => x"2025730a",
  1850 => x"00000000",
  1851 => x"20202020",
  1852 => x"20202020",
  1853 => x"73686f75",
  1854 => x"6c642062",
  1855 => x"653a2020",
  1856 => x"20444852",
  1857 => x"5953544f",
  1858 => x"4e452050",
  1859 => x"524f4752",
  1860 => x"414d2c20",
  1861 => x"534f4d45",
  1862 => x"20535452",
  1863 => x"494e470a",
  1864 => x"00000000",
  1865 => x"4e657874",
  1866 => x"5f507472",
  1867 => x"5f476c6f",
  1868 => x"622d3e0a",
  1869 => x"00000000",
  1870 => x"20202020",
  1871 => x"20202020",
  1872 => x"73686f75",
  1873 => x"6c642062",
  1874 => x"653a2020",
  1875 => x"2028696d",
  1876 => x"706c656d",
  1877 => x"656e7461",
  1878 => x"74696f6e",
  1879 => x"2d646570",
  1880 => x"656e6465",
  1881 => x"6e74292c",
  1882 => x"2073616d",
  1883 => x"65206173",
  1884 => x"2061626f",
  1885 => x"76650a00",
  1886 => x"496e745f",
  1887 => x"315f4c6f",
  1888 => x"633a2020",
  1889 => x"20202020",
  1890 => x"20202020",
  1891 => x"2025640a",
  1892 => x"00000000",
  1893 => x"496e745f",
  1894 => x"325f4c6f",
  1895 => x"633a2020",
  1896 => x"20202020",
  1897 => x"20202020",
  1898 => x"2025640a",
  1899 => x"00000000",
  1900 => x"496e745f",
  1901 => x"335f4c6f",
  1902 => x"633a2020",
  1903 => x"20202020",
  1904 => x"20202020",
  1905 => x"2025640a",
  1906 => x"00000000",
  1907 => x"456e756d",
  1908 => x"5f4c6f63",
  1909 => x"3a202020",
  1910 => x"20202020",
  1911 => x"20202020",
  1912 => x"2025640a",
  1913 => x"00000000",
  1914 => x"5374725f",
  1915 => x"315f4c6f",
  1916 => x"633a2020",
  1917 => x"20202020",
  1918 => x"20202020",
  1919 => x"2025730a",
  1920 => x"00000000",
  1921 => x"20202020",
  1922 => x"20202020",
  1923 => x"73686f75",
  1924 => x"6c642062",
  1925 => x"653a2020",
  1926 => x"20444852",
  1927 => x"5953544f",
  1928 => x"4e452050",
  1929 => x"524f4752",
  1930 => x"414d2c20",
  1931 => x"31275354",
  1932 => x"20535452",
  1933 => x"494e470a",
  1934 => x"00000000",
  1935 => x"5374725f",
  1936 => x"325f4c6f",
  1937 => x"633a2020",
  1938 => x"20202020",
  1939 => x"20202020",
  1940 => x"2025730a",
  1941 => x"00000000",
  1942 => x"20202020",
  1943 => x"20202020",
  1944 => x"73686f75",
  1945 => x"6c642062",
  1946 => x"653a2020",
  1947 => x"20444852",
  1948 => x"5953544f",
  1949 => x"4e452050",
  1950 => x"524f4752",
  1951 => x"414d2c20",
  1952 => x"32274e44",
  1953 => x"20535452",
  1954 => x"494e470a",
  1955 => x"00000000",
  1956 => x"55736572",
  1957 => x"2074696d",
  1958 => x"653a2025",
  1959 => x"640a0000",
  1960 => x"4d696372",
  1961 => x"6f736563",
  1962 => x"6f6e6473",
  1963 => x"20666f72",
  1964 => x"206f6e65",
  1965 => x"2072756e",
  1966 => x"20746872",
  1967 => x"6f756768",
  1968 => x"20446872",
  1969 => x"7973746f",
  1970 => x"6e653a20",
  1971 => x"00000000",
  1972 => x"2564200a",
  1973 => x"00000000",
  1974 => x"44687279",
  1975 => x"73746f6e",
  1976 => x"65732070",
  1977 => x"65722053",
  1978 => x"65636f6e",
  1979 => x"643a2020",
  1980 => x"20202020",
  1981 => x"20202020",
  1982 => x"20202020",
  1983 => x"20202020",
  1984 => x"20202020",
  1985 => x"00000000",
  1986 => x"56415820",
  1987 => x"4d495053",
  1988 => x"20726174",
  1989 => x"696e6720",
  1990 => x"2a203130",
  1991 => x"3030203d",
  1992 => x"20256420",
  1993 => x"0a000000",
  1994 => x"50726f67",
  1995 => x"72616d20",
  1996 => x"636f6d70",
  1997 => x"696c6564",
  1998 => x"20776974",
  1999 => x"686f7574",
  2000 => x"20277265",
  2001 => x"67697374",
  2002 => x"65722720",
  2003 => x"61747472",
  2004 => x"69627574",
  2005 => x"650a0000",
  2006 => x"4d656173",
  2007 => x"75726564",
  2008 => x"2074696d",
  2009 => x"6520746f",
  2010 => x"6f20736d",
  2011 => x"616c6c20",
  2012 => x"746f206f",
  2013 => x"62746169",
  2014 => x"6e206d65",
  2015 => x"616e696e",
  2016 => x"6766756c",
  2017 => x"20726573",
  2018 => x"756c7473",
  2019 => x"0a000000",
  2020 => x"506c6561",
  2021 => x"73652069",
  2022 => x"6e637265",
  2023 => x"61736520",
  2024 => x"6e756d62",
  2025 => x"6572206f",
  2026 => x"66207275",
  2027 => x"6e730a00",
  2028 => x"44485259",
  2029 => x"53544f4e",
  2030 => x"45205052",
  2031 => x"4f475241",
  2032 => x"4d2c2033",
  2033 => x"27524420",
  2034 => x"53545249",
  2035 => x"4e470000",
  2036 => x"30313233",
  2037 => x"34353637",
  2038 => x"38394142",
  2039 => x"43444546",
  2040 => x"00000000",
  2041 => x"64756d6d",
  2042 => x"792e6578",
  2043 => x"65000000",
  2044 => x"43000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"0000239c",
  2049 => x"000061a8",
  2050 => x"00000000",
  2051 => x"00001fe4",
  2052 => x"00002014",
  2053 => x"00000000",
  2054 => x"0000227c",
  2055 => x"000022d8",
  2056 => x"00002334",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00001ff0",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000001",
  2096 => x"330eabcd",
  2097 => x"1234e66d",
  2098 => x"deec0005",
  2099 => x"000b0000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000000",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"00000000",
  2209 => x"00000000",
  2210 => x"00000000",
  2211 => x"00000000",
  2212 => x"00000000",
  2213 => x"00000000",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"00000000",
  2217 => x"00000000",
  2218 => x"00000000",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000000",
  2244 => x"00000000",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"00000000",
  2262 => x"00000000",
  2263 => x"00000000",
  2264 => x"00000000",
  2265 => x"00000000",
  2266 => x"00000000",
  2267 => x"00000000",
  2268 => x"00000000",
  2269 => x"00000000",
  2270 => x"00000000",
  2271 => x"00000000",
  2272 => x"00000000",
  2273 => x"00000000",
  2274 => x"00000000",
  2275 => x"00000000",
  2276 => x"ffffffff",
  2277 => x"00000000",
  2278 => x"ffffffff",
  2279 => x"00000000",
  2280 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;


-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_ROM;

architecture arch of Dhrystone_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"80700b0b",
     2 => x"80c0fc0c",
     3 => x"3a0b0b0b",
     4 => x"a9cc0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"8f040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bb4",
   162 => x"d0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f7040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"df040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80c0f80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"83e13fac",
   257 => x"9d3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104b0",
   280 => x"08b408b8",
   281 => x"087575a3",
   282 => x"f22d5050",
   283 => x"b00856b8",
   284 => x"0cb40cb0",
   285 => x"0c5104b0",
   286 => x"08b408b8",
   287 => x"087575a2",
   288 => x"c02d5050",
   289 => x"b00856b8",
   290 => x"0cb40cb0",
   291 => x"0c5104b0",
   292 => x"08b408b8",
   293 => x"08aa932d",
   294 => x"b80cb40c",
   295 => x"b00c04fe",
   296 => x"3d0d0b0b",
   297 => x"80c8a808",
   298 => x"53841308",
   299 => x"70882a70",
   300 => x"81065152",
   301 => x"5270802e",
   302 => x"f0387181",
   303 => x"ff06b00c",
   304 => x"843d0d04",
   305 => x"ff3d0d0b",
   306 => x"0b80c8a8",
   307 => x"08527108",
   308 => x"70882a81",
   309 => x"32708106",
   310 => x"51515170",
   311 => x"f1387372",
   312 => x"0c833d0d",
   313 => x"0480c0f8",
   314 => x"08802ea4",
   315 => x"3880c0fc",
   316 => x"08822ebd",
   317 => x"38838080",
   318 => x"0b0b0b80",
   319 => x"c8a80c82",
   320 => x"a0800b80",
   321 => x"c8ac0c82",
   322 => x"90800b80",
   323 => x"c8b00c04",
   324 => x"f8808080",
   325 => x"a40b0b0b",
   326 => x"80c8a80c",
   327 => x"f8808082",
   328 => x"800b80c8",
   329 => x"ac0cf880",
   330 => x"8084800b",
   331 => x"80c8b00c",
   332 => x"0480c0a8",
   333 => x"808c0b0b",
   334 => x"0b80c8a8",
   335 => x"0c80c0a8",
   336 => x"80940b80",
   337 => x"c8ac0cb4",
   338 => x"e00b80c8",
   339 => x"b00c04f2",
   340 => x"3d0d6080",
   341 => x"c8ac0856",
   342 => x"5d82750c",
   343 => x"8059805a",
   344 => x"800b8f3d",
   345 => x"5d5b7a10",
   346 => x"10157008",
   347 => x"7108719f",
   348 => x"2c7e852b",
   349 => x"5855557d",
   350 => x"53595795",
   351 => x"cd3f7d7f",
   352 => x"7a72077c",
   353 => x"72077171",
   354 => x"60810541",
   355 => x"5f5d5b59",
   356 => x"5755817b",
   357 => x"278f3876",
   358 => x"7d0c7784",
   359 => x"1e0c7cb0",
   360 => x"0c903d0d",
   361 => x"0480c8ac",
   362 => x"0855ffba",
   363 => x"39ff3d0d",
   364 => x"80c8b433",
   365 => x"5170a738",
   366 => x"80c18408",
   367 => x"70085252",
   368 => x"70802e94",
   369 => x"38841280",
   370 => x"c1840c70",
   371 => x"2d80c184",
   372 => x"08700852",
   373 => x"5270ee38",
   374 => x"810b80c8",
   375 => x"b434833d",
   376 => x"0d040480",
   377 => x"3d0d0b0b",
   378 => x"80c8a408",
   379 => x"802e8e38",
   380 => x"0b0b0b0b",
   381 => x"800b802e",
   382 => x"09810685",
   383 => x"38823d0d",
   384 => x"040b0b80",
   385 => x"c8a4510b",
   386 => x"0b0bf3f4",
   387 => x"3f823d0d",
   388 => x"0404c008",
   389 => x"b00c0480",
   390 => x"3d0d80c1",
   391 => x"0b819898",
   392 => x"34800b81",
   393 => x"9ab00c70",
   394 => x"b00c823d",
   395 => x"0d04ff3d",
   396 => x"0d800b81",
   397 => x"98983352",
   398 => x"527080c1",
   399 => x"2e993871",
   400 => x"819ab008",
   401 => x"07819ab0",
   402 => x"0c80c20b",
   403 => x"81989c34",
   404 => x"70b00c83",
   405 => x"3d0d0481",
   406 => x"0b819ab0",
   407 => x"0807819a",
   408 => x"b00c80c2",
   409 => x"0b81989c",
   410 => x"3470b00c",
   411 => x"833d0d04",
   412 => x"fd3d0d75",
   413 => x"70088a05",
   414 => x"53538198",
   415 => x"98335170",
   416 => x"80c12e8b",
   417 => x"3873f338",
   418 => x"70b00c85",
   419 => x"3d0d04ff",
   420 => x"12708198",
   421 => x"94083174",
   422 => x"0cb00c85",
   423 => x"3d0d04fc",
   424 => x"3d0d8198",
   425 => x"c0085574",
   426 => x"802e8c38",
   427 => x"76750871",
   428 => x"0c8198c0",
   429 => x"0856548c",
   430 => x"15538198",
   431 => x"9408528a",
   432 => x"518cad3f",
   433 => x"73b00c86",
   434 => x"3d0d04fb",
   435 => x"3d0d7770",
   436 => x"085656b0",
   437 => x"538198c0",
   438 => x"08527451",
   439 => x"99c03f85",
   440 => x"0b8c170c",
   441 => x"850b8c16",
   442 => x"0c750875",
   443 => x"0c8198c0",
   444 => x"08547380",
   445 => x"2e8a3873",
   446 => x"08750c81",
   447 => x"98c00854",
   448 => x"8c145381",
   449 => x"98940852",
   450 => x"8a518be4",
   451 => x"3f841508",
   452 => x"ad38860b",
   453 => x"8c160c88",
   454 => x"15528816",
   455 => x"08518aea",
   456 => x"3f8198c0",
   457 => x"08700876",
   458 => x"0c548c15",
   459 => x"7054548a",
   460 => x"52730851",
   461 => x"8bba3f73",
   462 => x"b00c873d",
   463 => x"0d047508",
   464 => x"54b05373",
   465 => x"52755198",
   466 => x"d53f73b0",
   467 => x"0c873d0d",
   468 => x"04f33d0d",
   469 => x"88bd0bff",
   470 => x"880c8197",
   471 => x"ac0b8197",
   472 => x"e00c8197",
   473 => x"e40b8198",
   474 => x"c00c8197",
   475 => x"ac0b8197",
   476 => x"e40c800b",
   477 => x"8197e40b",
   478 => x"84050c82",
   479 => x"0b8197e4",
   480 => x"0b88050c",
   481 => x"a80b8197",
   482 => x"e40b8c05",
   483 => x"0c9f53b4",
   484 => x"e4528197",
   485 => x"f4519886",
   486 => x"3f9f53b5",
   487 => x"8452819a",
   488 => x"905197fa",
   489 => x"3f8a0b80",
   490 => x"d5f80cbf",
   491 => x"a8518ea5",
   492 => x"3fb5a451",
   493 => x"8e9f3fbf",
   494 => x"a8518e99",
   495 => x"3f80c18c",
   496 => x"08802e87",
   497 => x"d238b5d4",
   498 => x"518e8a3f",
   499 => x"bfa8518e",
   500 => x"843f80c1",
   501 => x"880852b6",
   502 => x"80518df9",
   503 => x"3fc00880",
   504 => x"c9980c81",
   505 => x"58800b80",
   506 => x"c1880825",
   507 => x"82d0388c",
   508 => x"3d5b80c1",
   509 => x"0b819898",
   510 => x"34810b81",
   511 => x"9ab00c80",
   512 => x"c20b8198",
   513 => x"9c34825c",
   514 => x"835a9f53",
   515 => x"b6b05281",
   516 => x"98a05197",
   517 => x"893f815d",
   518 => x"800b8198",
   519 => x"a053819a",
   520 => x"9052558b",
   521 => x"ae3fb008",
   522 => x"752e0981",
   523 => x"06833881",
   524 => x"5574819a",
   525 => x"b00c7b70",
   526 => x"57557483",
   527 => x"25a03874",
   528 => x"101015fd",
   529 => x"055e8f3d",
   530 => x"fc055383",
   531 => x"52755189",
   532 => x"9f3f811c",
   533 => x"705d7057",
   534 => x"55837524",
   535 => x"e2387d54",
   536 => x"745380c9",
   537 => x"9c528198",
   538 => x"c8518996",
   539 => x"3f8198c0",
   540 => x"08700857",
   541 => x"57b05376",
   542 => x"52755196",
   543 => x"a13f850b",
   544 => x"8c180c85",
   545 => x"0b8c170c",
   546 => x"7608760c",
   547 => x"8198c008",
   548 => x"5574802e",
   549 => x"8a387408",
   550 => x"760c8198",
   551 => x"c008558c",
   552 => x"15538198",
   553 => x"9408528a",
   554 => x"5188c53f",
   555 => x"84160887",
   556 => x"9038860b",
   557 => x"8c170c88",
   558 => x"16528817",
   559 => x"085187ca",
   560 => x"3f8198c0",
   561 => x"08700877",
   562 => x"0c558c16",
   563 => x"7054578a",
   564 => x"52760851",
   565 => x"889a3f80",
   566 => x"c10b8198",
   567 => x"9c335656",
   568 => x"757526a2",
   569 => x"3880c352",
   570 => x"755189ba",
   571 => x"3fb0087d",
   572 => x"2e86a038",
   573 => x"81167081",
   574 => x"ff068198",
   575 => x"9c335757",
   576 => x"57747627",
   577 => x"e038797c",
   578 => x"297e7072",
   579 => x"35705f72",
   580 => x"72317087",
   581 => x"29723153",
   582 => x"538a0581",
   583 => x"98983381",
   584 => x"9894085a",
   585 => x"5a525b55",
   586 => x"7680c12e",
   587 => x"86ab3878",
   588 => x"f7388118",
   589 => x"5880c188",
   590 => x"087825fd",
   591 => x"b538c008",
   592 => x"8197dc0c",
   593 => x"b6d0518b",
   594 => x"8c3fbfa8",
   595 => x"518b863f",
   596 => x"b6e0518b",
   597 => x"803fbfa8",
   598 => x"518afa3f",
   599 => x"81989408",
   600 => x"52b79851",
   601 => x"8aef3f85",
   602 => x"52b7b451",
   603 => x"8ae73f81",
   604 => x"9ab00852",
   605 => x"b7d0518a",
   606 => x"dc3f8152",
   607 => x"b7b4518a",
   608 => x"d43f8198",
   609 => x"983352b7",
   610 => x"ec518ac9",
   611 => x"3f80c152",
   612 => x"b888518a",
   613 => x"c03f8198",
   614 => x"9c3352b8",
   615 => x"a4518ab5",
   616 => x"3f80c252",
   617 => x"b888518a",
   618 => x"ac3f8198",
   619 => x"e80852b8",
   620 => x"c0518aa1",
   621 => x"3f8752b7",
   622 => x"b4518a99",
   623 => x"3f80d5f8",
   624 => x"0852b8dc",
   625 => x"518a8e3f",
   626 => x"b8f8518a",
   627 => x"883fb9a4",
   628 => x"518a823f",
   629 => x"8198c008",
   630 => x"70085357",
   631 => x"b9b05189",
   632 => x"f43fb9cc",
   633 => x"5189ee3f",
   634 => x"8198c008",
   635 => x"84110853",
   636 => x"5bba8051",
   637 => x"89df3f80",
   638 => x"52b7b451",
   639 => x"89d73f81",
   640 => x"98c00888",
   641 => x"11085358",
   642 => x"ba9c5189",
   643 => x"c83f8252",
   644 => x"b7b45189",
   645 => x"c03f8198",
   646 => x"c0088c11",
   647 => x"085359ba",
   648 => x"b85189b1",
   649 => x"3f9152b7",
   650 => x"b45189a9",
   651 => x"3f8198c0",
   652 => x"08900552",
   653 => x"bad45189",
   654 => x"9c3fbaf0",
   655 => x"5189963f",
   656 => x"bba85189",
   657 => x"903f8197",
   658 => x"e0087008",
   659 => x"5355b9b0",
   660 => x"5189823f",
   661 => x"bbbc5188",
   662 => x"fc3f8197",
   663 => x"e0088411",
   664 => x"085356ba",
   665 => x"805188ed",
   666 => x"3f8052b7",
   667 => x"b45188e5",
   668 => x"3f8197e0",
   669 => x"08881108",
   670 => x"5357ba9c",
   671 => x"5188d63f",
   672 => x"8152b7b4",
   673 => x"5188ce3f",
   674 => x"8197e008",
   675 => x"8c110853",
   676 => x"5bbab851",
   677 => x"88bf3f92",
   678 => x"52b7b451",
   679 => x"88b73f81",
   680 => x"97e00890",
   681 => x"0552bad4",
   682 => x"5188aa3f",
   683 => x"baf05188",
   684 => x"a43f7b52",
   685 => x"bbfc5188",
   686 => x"9c3f8552",
   687 => x"b7b45188",
   688 => x"943f7952",
   689 => x"bc985188",
   690 => x"8c3f8d52",
   691 => x"b7b45188",
   692 => x"843f7d52",
   693 => x"bcb45187",
   694 => x"fc3f8752",
   695 => x"b7b45187",
   696 => x"f43f7c52",
   697 => x"bcd05187",
   698 => x"ec3f8152",
   699 => x"b7b45187",
   700 => x"e43f819a",
   701 => x"9052bcec",
   702 => x"5187da3f",
   703 => x"bd885187",
   704 => x"d43f8198",
   705 => x"a052bdc0",
   706 => x"5187ca3f",
   707 => x"bddc5187",
   708 => x"c43fbfa8",
   709 => x"5187be3f",
   710 => x"8197dc08",
   711 => x"80c99808",
   712 => x"317080c9",
   713 => x"940c52be",
   714 => x"945187a9",
   715 => x"3f80c994",
   716 => x"085680f7",
   717 => x"762580e5",
   718 => x"3880c188",
   719 => x"08707787",
   720 => x"e8293580",
   721 => x"c98c0c76",
   722 => x"7187e829",
   723 => x"3580c990",
   724 => x"0c767184",
   725 => x"b9293581",
   726 => x"98c40c5a",
   727 => x"bea45186",
   728 => x"f43f80c9",
   729 => x"8c0852be",
   730 => x"d45186e9",
   731 => x"3fbedc51",
   732 => x"86e33f80",
   733 => x"c9900852",
   734 => x"bed45186",
   735 => x"d83f8198",
   736 => x"c40852bf",
   737 => x"8c5186cd",
   738 => x"3fbfa851",
   739 => x"86c73f80",
   740 => x"0bb00c8f",
   741 => x"3d0d04bf",
   742 => x"ac51f8ad",
   743 => x"39bfdc51",
   744 => x"86b33f80",
   745 => x"c0945186",
   746 => x"ac3fbfa8",
   747 => x"5186a63f",
   748 => x"80c99408",
   749 => x"80c18808",
   750 => x"707287e8",
   751 => x"293580c9",
   752 => x"8c0c7171",
   753 => x"87e82935",
   754 => x"80c9900c",
   755 => x"717184b9",
   756 => x"29358198",
   757 => x"c40c5b56",
   758 => x"bea45185",
   759 => x"f83f80c9",
   760 => x"8c0852be",
   761 => x"d45185ed",
   762 => x"3fbedc51",
   763 => x"85e73f80",
   764 => x"c9900852",
   765 => x"bed45185",
   766 => x"dc3f8198",
   767 => x"c40852bf",
   768 => x"8c5185d1",
   769 => x"3fbfa851",
   770 => x"85cb3f80",
   771 => x"0bb00c8f",
   772 => x"3d0d048f",
   773 => x"3df80552",
   774 => x"805180ee",
   775 => x"3f9f5380",
   776 => x"c0b45281",
   777 => x"98a0518e",
   778 => x"f53f7778",
   779 => x"8198940c",
   780 => x"81177081",
   781 => x"ff068198",
   782 => x"9c335858",
   783 => x"585af9c1",
   784 => x"39760856",
   785 => x"b0537552",
   786 => x"76518ed2",
   787 => x"3f80c10b",
   788 => x"81989c33",
   789 => x"5656f988",
   790 => x"39ff1570",
   791 => x"77317c0c",
   792 => x"59800b81",
   793 => x"19595980",
   794 => x"c1880878",
   795 => x"25f78338",
   796 => x"f9cc3902",
   797 => x"f8050d73",
   798 => x"82327030",
   799 => x"70720780",
   800 => x"25b00c52",
   801 => x"52028805",
   802 => x"0d0402f4",
   803 => x"050d7476",
   804 => x"71535452",
   805 => x"71822e83",
   806 => x"38835171",
   807 => x"812e9b38",
   808 => x"817226a0",
   809 => x"3871822e",
   810 => x"bc387184",
   811 => x"2eac3870",
   812 => x"730c70b0",
   813 => x"0c028c05",
   814 => x"0d0480e4",
   815 => x"0b819894",
   816 => x"08258c38",
   817 => x"80730c70",
   818 => x"b00c028c",
   819 => x"050d0483",
   820 => x"730c70b0",
   821 => x"0c028c05",
   822 => x"0d048273",
   823 => x"0c70b00c",
   824 => x"028c050d",
   825 => x"0481730c",
   826 => x"70b00c02",
   827 => x"8c050d04",
   828 => x"02fc050d",
   829 => x"74741482",
   830 => x"05710cb0",
   831 => x"0c028405",
   832 => x"0d0402d8",
   833 => x"050d7b7d",
   834 => x"7f618512",
   835 => x"70822b75",
   836 => x"11707471",
   837 => x"70840553",
   838 => x"0c5a5a5d",
   839 => x"5b760c79",
   840 => x"80f8180c",
   841 => x"79861252",
   842 => x"57585b59",
   843 => x"757725ac",
   844 => x"3881cc52",
   845 => x"7651a6bc",
   846 => x"2db0081a",
   847 => x"fc110881",
   848 => x"05fc120c",
   849 => x"79197008",
   850 => x"9fa0130c",
   851 => x"5b57850b",
   852 => x"8198940c",
   853 => x"76b00c02",
   854 => x"a8050d04",
   855 => x"b2527651",
   856 => x"a6bc2db0",
   857 => x"0817822b",
   858 => x"7a115153",
   859 => x"76737084",
   860 => x"05550c81",
   861 => x"14547574",
   862 => x"25f23881",
   863 => x"cc527651",
   864 => x"a6bc2db0",
   865 => x"081afc11",
   866 => x"088105fc",
   867 => x"120c7919",
   868 => x"70089fa0",
   869 => x"130c5b57",
   870 => x"850b8198",
   871 => x"940c76b0",
   872 => x"0c02a805",
   873 => x"0d0402f4",
   874 => x"050d0293",
   875 => x"05335180",
   876 => x"02840597",
   877 => x"05335452",
   878 => x"70732e89",
   879 => x"3871b00c",
   880 => x"028c050d",
   881 => x"04708198",
   882 => x"9834810b",
   883 => x"b00c028c",
   884 => x"050d0402",
   885 => x"dc050d7a",
   886 => x"7c595682",
   887 => x"0b831955",
   888 => x"55741670",
   889 => x"3375335b",
   890 => x"51537279",
   891 => x"2e80c738",
   892 => x"80c10b81",
   893 => x"16811656",
   894 => x"56578275",
   895 => x"25e338ff",
   896 => x"a9177081",
   897 => x"ff065559",
   898 => x"73822683",
   899 => x"38875581",
   900 => x"537680d2",
   901 => x"2e983877",
   902 => x"527551a8",
   903 => x"b72d8053",
   904 => x"72b00825",
   905 => x"89388715",
   906 => x"8198940c",
   907 => x"815372b0",
   908 => x"0c02a405",
   909 => x"0d047281",
   910 => x"98983482",
   911 => x"7525ffa1",
   912 => x"389bff04",
   913 => x"ff3d0d02",
   914 => x"8f053352",
   915 => x"ff840870",
   916 => x"882a7081",
   917 => x"06515151",
   918 => x"70802ef0",
   919 => x"3871ff84",
   920 => x"0c833d0d",
   921 => x"04fe3d0d",
   922 => x"74703352",
   923 => x"5370802e",
   924 => x"a1387052",
   925 => x"811353ff",
   926 => x"84087088",
   927 => x"2a708106",
   928 => x"51515170",
   929 => x"802ef038",
   930 => x"71ff840c",
   931 => x"72335271",
   932 => x"e338843d",
   933 => x"0d04ff3d",
   934 => x"0dff8408",
   935 => x"70892a70",
   936 => x"81065152",
   937 => x"5270802e",
   938 => x"f0387181",
   939 => x"ff06b00c",
   940 => x"833d0d04",
   941 => x"ff3d0d02",
   942 => x"8f053352",
   943 => x"ff840870",
   944 => x"882a7081",
   945 => x"06515151",
   946 => x"70802ef0",
   947 => x"3871ff84",
   948 => x"0c833d0d",
   949 => x"04f53d0d",
   950 => x"8e3d7070",
   951 => x"84055208",
   952 => x"9db45b55",
   953 => x"5b807470",
   954 => x"81055633",
   955 => x"755a5457",
   956 => x"72772ebe",
   957 => x"3872a52e",
   958 => x"09810680",
   959 => x"c5387770",
   960 => x"81055933",
   961 => x"537280e4",
   962 => x"2e81b638",
   963 => x"7280e424",
   964 => x"80c63872",
   965 => x"80e32ea1",
   966 => x"388052a5",
   967 => x"51782d80",
   968 => x"52725178",
   969 => x"2d821757",
   970 => x"77708105",
   971 => x"59335372",
   972 => x"c43876b0",
   973 => x"0c8d3d0d",
   974 => x"047a841c",
   975 => x"83123355",
   976 => x"5c568052",
   977 => x"7251782d",
   978 => x"81177870",
   979 => x"81055a33",
   980 => x"545772ff",
   981 => x"a038db39",
   982 => x"7280f32e",
   983 => x"098106ff",
   984 => x"b8387a84",
   985 => x"1c710858",
   986 => x"5c548076",
   987 => x"335b5579",
   988 => x"752e8d38",
   989 => x"81157017",
   990 => x"7033555b",
   991 => x"5572f538",
   992 => x"ff155480",
   993 => x"7525ffa0",
   994 => x"38757081",
   995 => x"05573353",
   996 => x"80527251",
   997 => x"782d8117",
   998 => x"74ff1656",
   999 => x"56578075",
  1000 => x"25ff8538",
  1001 => x"75708105",
  1002 => x"57335380",
  1003 => x"52725178",
  1004 => x"2d811774",
  1005 => x"ff165656",
  1006 => x"57748024",
  1007 => x"cc38fee8",
  1008 => x"397a841c",
  1009 => x"7108819a",
  1010 => x"c40b80c8",
  1011 => x"b8545d56",
  1012 => x"5c558056",
  1013 => x"73762e09",
  1014 => x"8106b838",
  1015 => x"b00b80c8",
  1016 => x"b8348115",
  1017 => x"55ff1555",
  1018 => x"74337a70",
  1019 => x"81055c34",
  1020 => x"81165674",
  1021 => x"80c8b82e",
  1022 => x"098106e9",
  1023 => x"38807a34",
  1024 => x"75819ac4",
  1025 => x"0bff1256",
  1026 => x"57557480",
  1027 => x"24fefa38",
  1028 => x"fe963973",
  1029 => x"8f0680c0",
  1030 => x"d4055372",
  1031 => x"33757081",
  1032 => x"05573473",
  1033 => x"842a5473",
  1034 => x"ea387480",
  1035 => x"c8b82ecd",
  1036 => x"38ff1555",
  1037 => x"74337a70",
  1038 => x"81055c34",
  1039 => x"81165674",
  1040 => x"80c8b82e",
  1041 => x"ffb738ff",
  1042 => x"9c39bc08",
  1043 => x"02bc0cf5",
  1044 => x"3d0dbc08",
  1045 => x"9405089d",
  1046 => x"38bc088c",
  1047 => x"0508bc08",
  1048 => x"900508bc",
  1049 => x"08880508",
  1050 => x"58565473",
  1051 => x"760c7484",
  1052 => x"170c81bf",
  1053 => x"39800bbc",
  1054 => x"08f0050c",
  1055 => x"800bbc08",
  1056 => x"f4050cbc",
  1057 => x"088c0508",
  1058 => x"bc089005",
  1059 => x"08565473",
  1060 => x"bc08f005",
  1061 => x"0c74bc08",
  1062 => x"f4050cbc",
  1063 => x"08f805bc",
  1064 => x"08f00556",
  1065 => x"56887054",
  1066 => x"75537652",
  1067 => x"5485ef3f",
  1068 => x"a00bbc08",
  1069 => x"94050831",
  1070 => x"bc08ec05",
  1071 => x"0cbc08ec",
  1072 => x"05088024",
  1073 => x"9d38800b",
  1074 => x"bc08f405",
  1075 => x"0cbc08ec",
  1076 => x"050830bc",
  1077 => x"08fc0508",
  1078 => x"712bbc08",
  1079 => x"f0050c54",
  1080 => x"b939bc08",
  1081 => x"fc0508bc",
  1082 => x"08ec0508",
  1083 => x"2abc08e8",
  1084 => x"050cbc08",
  1085 => x"fc0508bc",
  1086 => x"08940508",
  1087 => x"2bbc08f4",
  1088 => x"050cbc08",
  1089 => x"f80508bc",
  1090 => x"08940508",
  1091 => x"2b70bc08",
  1092 => x"e8050807",
  1093 => x"bc08f005",
  1094 => x"0c54bc08",
  1095 => x"f00508bc",
  1096 => x"08f40508",
  1097 => x"bc088805",
  1098 => x"08585654",
  1099 => x"73760c74",
  1100 => x"84170cbc",
  1101 => x"08880508",
  1102 => x"b00c8d3d",
  1103 => x"0dbc0c04",
  1104 => x"bc0802bc",
  1105 => x"0cf93d0d",
  1106 => x"800bbc08",
  1107 => x"fc050cbc",
  1108 => x"08880508",
  1109 => x"8025ab38",
  1110 => x"bc088805",
  1111 => x"0830bc08",
  1112 => x"88050c80",
  1113 => x"0bbc08f4",
  1114 => x"050cbc08",
  1115 => x"fc050888",
  1116 => x"38810bbc",
  1117 => x"08f4050c",
  1118 => x"bc08f405",
  1119 => x"08bc08fc",
  1120 => x"050cbc08",
  1121 => x"8c050880",
  1122 => x"25ab38bc",
  1123 => x"088c0508",
  1124 => x"30bc088c",
  1125 => x"050c800b",
  1126 => x"bc08f005",
  1127 => x"0cbc08fc",
  1128 => x"05088838",
  1129 => x"810bbc08",
  1130 => x"f0050cbc",
  1131 => x"08f00508",
  1132 => x"bc08fc05",
  1133 => x"0c8053bc",
  1134 => x"088c0508",
  1135 => x"52bc0888",
  1136 => x"05085181",
  1137 => x"a73fb008",
  1138 => x"70bc08f8",
  1139 => x"050c54bc",
  1140 => x"08fc0508",
  1141 => x"802e8c38",
  1142 => x"bc08f805",
  1143 => x"0830bc08",
  1144 => x"f8050cbc",
  1145 => x"08f80508",
  1146 => x"70b00c54",
  1147 => x"893d0dbc",
  1148 => x"0c04bc08",
  1149 => x"02bc0cfb",
  1150 => x"3d0d800b",
  1151 => x"bc08fc05",
  1152 => x"0cbc0888",
  1153 => x"05088025",
  1154 => x"9338bc08",
  1155 => x"88050830",
  1156 => x"bc088805",
  1157 => x"0c810bbc",
  1158 => x"08fc050c",
  1159 => x"bc088c05",
  1160 => x"0880258c",
  1161 => x"38bc088c",
  1162 => x"050830bc",
  1163 => x"088c050c",
  1164 => x"8153bc08",
  1165 => x"8c050852",
  1166 => x"bc088805",
  1167 => x"0851ad3f",
  1168 => x"b00870bc",
  1169 => x"08f8050c",
  1170 => x"54bc08fc",
  1171 => x"0508802e",
  1172 => x"8c38bc08",
  1173 => x"f8050830",
  1174 => x"bc08f805",
  1175 => x"0cbc08f8",
  1176 => x"050870b0",
  1177 => x"0c54873d",
  1178 => x"0dbc0c04",
  1179 => x"bc0802bc",
  1180 => x"0cfd3d0d",
  1181 => x"810bbc08",
  1182 => x"fc050c80",
  1183 => x"0bbc08f8",
  1184 => x"050cbc08",
  1185 => x"8c0508bc",
  1186 => x"08880508",
  1187 => x"27ac38bc",
  1188 => x"08fc0508",
  1189 => x"802ea338",
  1190 => x"800bbc08",
  1191 => x"8c050824",
  1192 => x"9938bc08",
  1193 => x"8c050810",
  1194 => x"bc088c05",
  1195 => x"0cbc08fc",
  1196 => x"050810bc",
  1197 => x"08fc050c",
  1198 => x"c939bc08",
  1199 => x"fc050880",
  1200 => x"2e80c938",
  1201 => x"bc088c05",
  1202 => x"08bc0888",
  1203 => x"050826a1",
  1204 => x"38bc0888",
  1205 => x"0508bc08",
  1206 => x"8c050831",
  1207 => x"bc088805",
  1208 => x"0cbc08f8",
  1209 => x"0508bc08",
  1210 => x"fc050807",
  1211 => x"bc08f805",
  1212 => x"0cbc08fc",
  1213 => x"0508812a",
  1214 => x"bc08fc05",
  1215 => x"0cbc088c",
  1216 => x"0508812a",
  1217 => x"bc088c05",
  1218 => x"0cffaf39",
  1219 => x"bc089005",
  1220 => x"08802e8f",
  1221 => x"38bc0888",
  1222 => x"050870bc",
  1223 => x"08f4050c",
  1224 => x"518d39bc",
  1225 => x"08f80508",
  1226 => x"70bc08f4",
  1227 => x"050c51bc",
  1228 => x"08f40508",
  1229 => x"b00c853d",
  1230 => x"0dbc0c04",
  1231 => x"bc0802bc",
  1232 => x"0cff3d0d",
  1233 => x"800bbc08",
  1234 => x"fc050cbc",
  1235 => x"08880508",
  1236 => x"8106ff11",
  1237 => x"700970bc",
  1238 => x"088c0508",
  1239 => x"06bc08fc",
  1240 => x"050811bc",
  1241 => x"08fc050c",
  1242 => x"bc088805",
  1243 => x"08812abc",
  1244 => x"0888050c",
  1245 => x"bc088c05",
  1246 => x"0810bc08",
  1247 => x"8c050c51",
  1248 => x"515151bc",
  1249 => x"08880508",
  1250 => x"802e8438",
  1251 => x"ffbd39bc",
  1252 => x"08fc0508",
  1253 => x"70b00c51",
  1254 => x"833d0dbc",
  1255 => x"0c04fc3d",
  1256 => x"0d767079",
  1257 => x"7b555555",
  1258 => x"558f7227",
  1259 => x"8c387275",
  1260 => x"07830651",
  1261 => x"70802ea7",
  1262 => x"38ff1252",
  1263 => x"71ff2e98",
  1264 => x"38727081",
  1265 => x"05543374",
  1266 => x"70810556",
  1267 => x"34ff1252",
  1268 => x"71ff2e09",
  1269 => x"8106ea38",
  1270 => x"74b00c86",
  1271 => x"3d0d0474",
  1272 => x"51727084",
  1273 => x"05540871",
  1274 => x"70840553",
  1275 => x"0c727084",
  1276 => x"05540871",
  1277 => x"70840553",
  1278 => x"0c727084",
  1279 => x"05540871",
  1280 => x"70840553",
  1281 => x"0c727084",
  1282 => x"05540871",
  1283 => x"70840553",
  1284 => x"0cf01252",
  1285 => x"718f26c9",
  1286 => x"38837227",
  1287 => x"95387270",
  1288 => x"84055408",
  1289 => x"71708405",
  1290 => x"530cfc12",
  1291 => x"52718326",
  1292 => x"ed387054",
  1293 => x"ff8339fb",
  1294 => x"3d0d7779",
  1295 => x"70720783",
  1296 => x"06535452",
  1297 => x"70933871",
  1298 => x"73730854",
  1299 => x"56547173",
  1300 => x"082e80c4",
  1301 => x"38737554",
  1302 => x"52713370",
  1303 => x"81ff0652",
  1304 => x"5470802e",
  1305 => x"9d387233",
  1306 => x"5570752e",
  1307 => x"09810695",
  1308 => x"38811281",
  1309 => x"14713370",
  1310 => x"81ff0654",
  1311 => x"56545270",
  1312 => x"e5387233",
  1313 => x"557381ff",
  1314 => x"067581ff",
  1315 => x"06717131",
  1316 => x"b00c5252",
  1317 => x"873d0d04",
  1318 => x"710970f7",
  1319 => x"fbfdff14",
  1320 => x"0670f884",
  1321 => x"82818006",
  1322 => x"51515170",
  1323 => x"97388414",
  1324 => x"84167108",
  1325 => x"54565471",
  1326 => x"75082edc",
  1327 => x"38737554",
  1328 => x"52ff9639",
  1329 => x"800bb00c",
  1330 => x"873d0d04",
  1331 => x"fd3d0d80",
  1332 => x"0b80c0fc",
  1333 => x"08545472",
  1334 => x"812e9b38",
  1335 => x"7380c988",
  1336 => x"0ce0823f",
  1337 => x"de9a3f80",
  1338 => x"c1905281",
  1339 => x"51e4e23f",
  1340 => x"b0085187",
  1341 => x"9b3f7280",
  1342 => x"c9880cdf",
  1343 => x"e83fde80",
  1344 => x"3f80c190",
  1345 => x"528151e4",
  1346 => x"c83fb008",
  1347 => x"5187813f",
  1348 => x"00ff3900",
  1349 => x"ff39f53d",
  1350 => x"0d7e6080",
  1351 => x"c9880870",
  1352 => x"5b585b5b",
  1353 => x"7580c238",
  1354 => x"777a25a1",
  1355 => x"38771b70",
  1356 => x"337081ff",
  1357 => x"06585859",
  1358 => x"758a2e98",
  1359 => x"387681ff",
  1360 => x"0651df80",
  1361 => x"3f811858",
  1362 => x"797824e1",
  1363 => x"3879b00c",
  1364 => x"8d3d0d04",
  1365 => x"8d51deec",
  1366 => x"3f783370",
  1367 => x"81ff0652",
  1368 => x"57dee13f",
  1369 => x"811858e0",
  1370 => x"3979557a",
  1371 => x"547d5385",
  1372 => x"528d3dfc",
  1373 => x"0551ddc9",
  1374 => x"3fb00856",
  1375 => x"868b3f7b",
  1376 => x"b0080c75",
  1377 => x"b00c8d3d",
  1378 => x"0d04f63d",
  1379 => x"0d7d7f80",
  1380 => x"c9880870",
  1381 => x"5b585a5a",
  1382 => x"7580c138",
  1383 => x"777925b3",
  1384 => x"38ddfc3f",
  1385 => x"b00881ff",
  1386 => x"06708d32",
  1387 => x"7030709f",
  1388 => x"2a515157",
  1389 => x"57768a2e",
  1390 => x"80c33875",
  1391 => x"802ebe38",
  1392 => x"771a5676",
  1393 => x"76347651",
  1394 => x"ddfa3f81",
  1395 => x"18587878",
  1396 => x"24cf3877",
  1397 => x"5675b00c",
  1398 => x"8c3d0d04",
  1399 => x"78557954",
  1400 => x"7c538452",
  1401 => x"8c3dfc05",
  1402 => x"51dcd63f",
  1403 => x"b0085685",
  1404 => x"983f7ab0",
  1405 => x"080c75b0",
  1406 => x"0c8c3d0d",
  1407 => x"04771a56",
  1408 => x"8a763481",
  1409 => x"18588d51",
  1410 => x"ddba3f8a",
  1411 => x"51ddb53f",
  1412 => x"7756c239",
  1413 => x"f93d0d79",
  1414 => x"5780c988",
  1415 => x"08802eac",
  1416 => x"38765187",
  1417 => x"9e3f7b56",
  1418 => x"7a55b008",
  1419 => x"81055476",
  1420 => x"53825289",
  1421 => x"3dfc0551",
  1422 => x"dc873fb0",
  1423 => x"085784c9",
  1424 => x"3f77b008",
  1425 => x"0c76b00c",
  1426 => x"893d0d04",
  1427 => x"84bb3f85",
  1428 => x"0bb0080c",
  1429 => x"ff0bb00c",
  1430 => x"893d0d04",
  1431 => x"fb3d0d80",
  1432 => x"c9880870",
  1433 => x"56547388",
  1434 => x"3874b00c",
  1435 => x"873d0d04",
  1436 => x"77538352",
  1437 => x"873dfc05",
  1438 => x"51dbc63f",
  1439 => x"b0085484",
  1440 => x"883f75b0",
  1441 => x"080c73b0",
  1442 => x"0c873d0d",
  1443 => x"04ff0bb0",
  1444 => x"0c04fb3d",
  1445 => x"0d775580",
  1446 => x"c9880880",
  1447 => x"2ea83874",
  1448 => x"5186a03f",
  1449 => x"b0088105",
  1450 => x"54745387",
  1451 => x"52873dfc",
  1452 => x"0551db8d",
  1453 => x"3fb00855",
  1454 => x"83cf3f75",
  1455 => x"b0080c74",
  1456 => x"b00c873d",
  1457 => x"0d0483c1",
  1458 => x"3f850bb0",
  1459 => x"080cff0b",
  1460 => x"b00c873d",
  1461 => x"0d04fa3d",
  1462 => x"0d80c988",
  1463 => x"08802ea2",
  1464 => x"387a5579",
  1465 => x"54785386",
  1466 => x"52883dfc",
  1467 => x"0551dad1",
  1468 => x"3fb00856",
  1469 => x"83933f76",
  1470 => x"b0080c75",
  1471 => x"b00c883d",
  1472 => x"0d048385",
  1473 => x"3f9d0bb0",
  1474 => x"080cff0b",
  1475 => x"b00c883d",
  1476 => x"0d04fb3d",
  1477 => x"0d777956",
  1478 => x"56807054",
  1479 => x"54737525",
  1480 => x"9f387410",
  1481 => x"1010f805",
  1482 => x"52721670",
  1483 => x"3370742b",
  1484 => x"76078116",
  1485 => x"f8165656",
  1486 => x"56515174",
  1487 => x"7324ea38",
  1488 => x"73b00c87",
  1489 => x"3d0d04fc",
  1490 => x"3d0d7678",
  1491 => x"5555bc53",
  1492 => x"80527351",
  1493 => x"83de3f84",
  1494 => x"527451ff",
  1495 => x"b53fb008",
  1496 => x"74238452",
  1497 => x"841551ff",
  1498 => x"a93fb008",
  1499 => x"82152384",
  1500 => x"52881551",
  1501 => x"ff9c3fb0",
  1502 => x"0884150c",
  1503 => x"84528c15",
  1504 => x"51ff8f3f",
  1505 => x"b0088815",
  1506 => x"23845290",
  1507 => x"1551ff82",
  1508 => x"3fb0088a",
  1509 => x"15238452",
  1510 => x"941551fe",
  1511 => x"f53fb008",
  1512 => x"8c152384",
  1513 => x"52981551",
  1514 => x"fee83fb0",
  1515 => x"088e1523",
  1516 => x"88529c15",
  1517 => x"51fedb3f",
  1518 => x"b0089015",
  1519 => x"0c863d0d",
  1520 => x"04e93d0d",
  1521 => x"6a80c988",
  1522 => x"08575775",
  1523 => x"933880c0",
  1524 => x"800b8418",
  1525 => x"0c75ac18",
  1526 => x"0c75b00c",
  1527 => x"993d0d04",
  1528 => x"893d7055",
  1529 => x"6a54558a",
  1530 => x"52993dff",
  1531 => x"bc0551d8",
  1532 => x"d03fb008",
  1533 => x"77537552",
  1534 => x"56fecc3f",
  1535 => x"818b3f77",
  1536 => x"b0080c75",
  1537 => x"b00c993d",
  1538 => x"0d04e93d",
  1539 => x"0d695780",
  1540 => x"c9880880",
  1541 => x"2eb53876",
  1542 => x"5183a83f",
  1543 => x"893d7056",
  1544 => x"b0088105",
  1545 => x"55775456",
  1546 => x"8f52993d",
  1547 => x"ffbc0551",
  1548 => x"d88f3fb0",
  1549 => x"086b5376",
  1550 => x"5257fe8b",
  1551 => x"3f80ca3f",
  1552 => x"77b0080c",
  1553 => x"76b00c99",
  1554 => x"3d0d04bd",
  1555 => x"3f850bb0",
  1556 => x"080cff0b",
  1557 => x"b00c993d",
  1558 => x"0d04fc3d",
  1559 => x"0d815480",
  1560 => x"c9880888",
  1561 => x"3873b00c",
  1562 => x"863d0d04",
  1563 => x"765397b9",
  1564 => x"52863dfc",
  1565 => x"0551d7c9",
  1566 => x"3fb00854",
  1567 => x"8c3f74b0",
  1568 => x"080c73b0",
  1569 => x"0c863d0d",
  1570 => x"0480c194",
  1571 => x"08b00c04",
  1572 => x"f73d0d7b",
  1573 => x"80c19408",
  1574 => x"82c81108",
  1575 => x"5a545a77",
  1576 => x"802e80da",
  1577 => x"38818818",
  1578 => x"841908ff",
  1579 => x"0581712b",
  1580 => x"59555980",
  1581 => x"742480ea",
  1582 => x"38807424",
  1583 => x"b5387382",
  1584 => x"2b781188",
  1585 => x"05565681",
  1586 => x"80190877",
  1587 => x"06537280",
  1588 => x"2eb63878",
  1589 => x"16700853",
  1590 => x"53795174",
  1591 => x"0853722d",
  1592 => x"ff14fc17",
  1593 => x"fc177981",
  1594 => x"2c5a5757",
  1595 => x"54738025",
  1596 => x"d6387708",
  1597 => x"5877ffad",
  1598 => x"3880c194",
  1599 => x"0853bc13",
  1600 => x"08a53879",
  1601 => x"51f8893f",
  1602 => x"74085372",
  1603 => x"2dff14fc",
  1604 => x"17fc1779",
  1605 => x"812c5a57",
  1606 => x"57547380",
  1607 => x"25ffa838",
  1608 => x"d1398057",
  1609 => x"ff933972",
  1610 => x"51bc1308",
  1611 => x"53722d79",
  1612 => x"51f7dd3f",
  1613 => x"fc3d0d76",
  1614 => x"7971028c",
  1615 => x"059f0533",
  1616 => x"57555355",
  1617 => x"8372278a",
  1618 => x"38748306",
  1619 => x"5170802e",
  1620 => x"a238ff12",
  1621 => x"5271ff2e",
  1622 => x"93387373",
  1623 => x"70810555",
  1624 => x"34ff1252",
  1625 => x"71ff2e09",
  1626 => x"8106ef38",
  1627 => x"74b00c86",
  1628 => x"3d0d0474",
  1629 => x"74882b75",
  1630 => x"07707190",
  1631 => x"2b075154",
  1632 => x"518f7227",
  1633 => x"a5387271",
  1634 => x"70840553",
  1635 => x"0c727170",
  1636 => x"8405530c",
  1637 => x"72717084",
  1638 => x"05530c72",
  1639 => x"71708405",
  1640 => x"530cf012",
  1641 => x"52718f26",
  1642 => x"dd388372",
  1643 => x"27903872",
  1644 => x"71708405",
  1645 => x"530cfc12",
  1646 => x"52718326",
  1647 => x"f2387053",
  1648 => x"ff9039fd",
  1649 => x"3d0d7570",
  1650 => x"71830653",
  1651 => x"555270b8",
  1652 => x"38717008",
  1653 => x"7009f7fb",
  1654 => x"fdff1206",
  1655 => x"70f88482",
  1656 => x"81800651",
  1657 => x"51525370",
  1658 => x"9d388413",
  1659 => x"70087009",
  1660 => x"f7fbfdff",
  1661 => x"120670f8",
  1662 => x"84828180",
  1663 => x"06515152",
  1664 => x"5370802e",
  1665 => x"e5387252",
  1666 => x"71335170",
  1667 => x"802e8a38",
  1668 => x"81127033",
  1669 => x"525270f8",
  1670 => x"38717431",
  1671 => x"b00c853d",
  1672 => x"0d04ff3d",
  1673 => x"0d80c898",
  1674 => x"0bfc0570",
  1675 => x"08525270",
  1676 => x"ff2e9138",
  1677 => x"702dfc12",
  1678 => x"70085252",
  1679 => x"70ff2e09",
  1680 => x"8106f138",
  1681 => x"833d0d04",
  1682 => x"04d6e23f",
  1683 => x"04000000",
  1684 => x"00ffffff",
  1685 => x"ff00ffff",
  1686 => x"ffff00ff",
  1687 => x"ffffff00",
  1688 => x"00000040",
  1689 => x"44485259",
  1690 => x"53544f4e",
  1691 => x"45205052",
  1692 => x"4f475241",
  1693 => x"4d2c2053",
  1694 => x"4f4d4520",
  1695 => x"53545249",
  1696 => x"4e470000",
  1697 => x"44485259",
  1698 => x"53544f4e",
  1699 => x"45205052",
  1700 => x"4f475241",
  1701 => x"4d2c2031",
  1702 => x"27535420",
  1703 => x"53545249",
  1704 => x"4e470000",
  1705 => x"44687279",
  1706 => x"73746f6e",
  1707 => x"65204265",
  1708 => x"6e63686d",
  1709 => x"61726b2c",
  1710 => x"20566572",
  1711 => x"73696f6e",
  1712 => x"20322e31",
  1713 => x"20284c61",
  1714 => x"6e677561",
  1715 => x"67653a20",
  1716 => x"43290a00",
  1717 => x"50726f67",
  1718 => x"72616d20",
  1719 => x"636f6d70",
  1720 => x"696c6564",
  1721 => x"20776974",
  1722 => x"68202772",
  1723 => x"65676973",
  1724 => x"74657227",
  1725 => x"20617474",
  1726 => x"72696275",
  1727 => x"74650a00",
  1728 => x"45786563",
  1729 => x"7574696f",
  1730 => x"6e207374",
  1731 => x"61727473",
  1732 => x"2c202564",
  1733 => x"2072756e",
  1734 => x"73207468",
  1735 => x"726f7567",
  1736 => x"68204468",
  1737 => x"72797374",
  1738 => x"6f6e650a",
  1739 => x"00000000",
  1740 => x"44485259",
  1741 => x"53544f4e",
  1742 => x"45205052",
  1743 => x"4f475241",
  1744 => x"4d2c2032",
  1745 => x"274e4420",
  1746 => x"53545249",
  1747 => x"4e470000",
  1748 => x"45786563",
  1749 => x"7574696f",
  1750 => x"6e20656e",
  1751 => x"64730a00",
  1752 => x"46696e61",
  1753 => x"6c207661",
  1754 => x"6c756573",
  1755 => x"206f6620",
  1756 => x"74686520",
  1757 => x"76617269",
  1758 => x"61626c65",
  1759 => x"73207573",
  1760 => x"65642069",
  1761 => x"6e207468",
  1762 => x"65206265",
  1763 => x"6e63686d",
  1764 => x"61726b3a",
  1765 => x"0a000000",
  1766 => x"496e745f",
  1767 => x"476c6f62",
  1768 => x"3a202020",
  1769 => x"20202020",
  1770 => x"20202020",
  1771 => x"2025640a",
  1772 => x"00000000",
  1773 => x"20202020",
  1774 => x"20202020",
  1775 => x"73686f75",
  1776 => x"6c642062",
  1777 => x"653a2020",
  1778 => x"2025640a",
  1779 => x"00000000",
  1780 => x"426f6f6c",
  1781 => x"5f476c6f",
  1782 => x"623a2020",
  1783 => x"20202020",
  1784 => x"20202020",
  1785 => x"2025640a",
  1786 => x"00000000",
  1787 => x"43685f31",
  1788 => x"5f476c6f",
  1789 => x"623a2020",
  1790 => x"20202020",
  1791 => x"20202020",
  1792 => x"2025630a",
  1793 => x"00000000",
  1794 => x"20202020",
  1795 => x"20202020",
  1796 => x"73686f75",
  1797 => x"6c642062",
  1798 => x"653a2020",
  1799 => x"2025630a",
  1800 => x"00000000",
  1801 => x"43685f32",
  1802 => x"5f476c6f",
  1803 => x"623a2020",
  1804 => x"20202020",
  1805 => x"20202020",
  1806 => x"2025630a",
  1807 => x"00000000",
  1808 => x"4172725f",
  1809 => x"315f476c",
  1810 => x"6f625b38",
  1811 => x"5d3a2020",
  1812 => x"20202020",
  1813 => x"2025640a",
  1814 => x"00000000",
  1815 => x"4172725f",
  1816 => x"325f476c",
  1817 => x"6f625b38",
  1818 => x"5d5b375d",
  1819 => x"3a202020",
  1820 => x"2025640a",
  1821 => x"00000000",
  1822 => x"20202020",
  1823 => x"20202020",
  1824 => x"73686f75",
  1825 => x"6c642062",
  1826 => x"653a2020",
  1827 => x"204e756d",
  1828 => x"6265725f",
  1829 => x"4f665f52",
  1830 => x"756e7320",
  1831 => x"2b203130",
  1832 => x"0a000000",
  1833 => x"5074725f",
  1834 => x"476c6f62",
  1835 => x"2d3e0a00",
  1836 => x"20205074",
  1837 => x"725f436f",
  1838 => x"6d703a20",
  1839 => x"20202020",
  1840 => x"20202020",
  1841 => x"2025640a",
  1842 => x"00000000",
  1843 => x"20202020",
  1844 => x"20202020",
  1845 => x"73686f75",
  1846 => x"6c642062",
  1847 => x"653a2020",
  1848 => x"2028696d",
  1849 => x"706c656d",
  1850 => x"656e7461",
  1851 => x"74696f6e",
  1852 => x"2d646570",
  1853 => x"656e6465",
  1854 => x"6e74290a",
  1855 => x"00000000",
  1856 => x"20204469",
  1857 => x"7363723a",
  1858 => x"20202020",
  1859 => x"20202020",
  1860 => x"20202020",
  1861 => x"2025640a",
  1862 => x"00000000",
  1863 => x"2020456e",
  1864 => x"756d5f43",
  1865 => x"6f6d703a",
  1866 => x"20202020",
  1867 => x"20202020",
  1868 => x"2025640a",
  1869 => x"00000000",
  1870 => x"2020496e",
  1871 => x"745f436f",
  1872 => x"6d703a20",
  1873 => x"20202020",
  1874 => x"20202020",
  1875 => x"2025640a",
  1876 => x"00000000",
  1877 => x"20205374",
  1878 => x"725f436f",
  1879 => x"6d703a20",
  1880 => x"20202020",
  1881 => x"20202020",
  1882 => x"2025730a",
  1883 => x"00000000",
  1884 => x"20202020",
  1885 => x"20202020",
  1886 => x"73686f75",
  1887 => x"6c642062",
  1888 => x"653a2020",
  1889 => x"20444852",
  1890 => x"5953544f",
  1891 => x"4e452050",
  1892 => x"524f4752",
  1893 => x"414d2c20",
  1894 => x"534f4d45",
  1895 => x"20535452",
  1896 => x"494e470a",
  1897 => x"00000000",
  1898 => x"4e657874",
  1899 => x"5f507472",
  1900 => x"5f476c6f",
  1901 => x"622d3e0a",
  1902 => x"00000000",
  1903 => x"20202020",
  1904 => x"20202020",
  1905 => x"73686f75",
  1906 => x"6c642062",
  1907 => x"653a2020",
  1908 => x"2028696d",
  1909 => x"706c656d",
  1910 => x"656e7461",
  1911 => x"74696f6e",
  1912 => x"2d646570",
  1913 => x"656e6465",
  1914 => x"6e74292c",
  1915 => x"2073616d",
  1916 => x"65206173",
  1917 => x"2061626f",
  1918 => x"76650a00",
  1919 => x"496e745f",
  1920 => x"315f4c6f",
  1921 => x"633a2020",
  1922 => x"20202020",
  1923 => x"20202020",
  1924 => x"2025640a",
  1925 => x"00000000",
  1926 => x"496e745f",
  1927 => x"325f4c6f",
  1928 => x"633a2020",
  1929 => x"20202020",
  1930 => x"20202020",
  1931 => x"2025640a",
  1932 => x"00000000",
  1933 => x"496e745f",
  1934 => x"335f4c6f",
  1935 => x"633a2020",
  1936 => x"20202020",
  1937 => x"20202020",
  1938 => x"2025640a",
  1939 => x"00000000",
  1940 => x"456e756d",
  1941 => x"5f4c6f63",
  1942 => x"3a202020",
  1943 => x"20202020",
  1944 => x"20202020",
  1945 => x"2025640a",
  1946 => x"00000000",
  1947 => x"5374725f",
  1948 => x"315f4c6f",
  1949 => x"633a2020",
  1950 => x"20202020",
  1951 => x"20202020",
  1952 => x"2025730a",
  1953 => x"00000000",
  1954 => x"20202020",
  1955 => x"20202020",
  1956 => x"73686f75",
  1957 => x"6c642062",
  1958 => x"653a2020",
  1959 => x"20444852",
  1960 => x"5953544f",
  1961 => x"4e452050",
  1962 => x"524f4752",
  1963 => x"414d2c20",
  1964 => x"31275354",
  1965 => x"20535452",
  1966 => x"494e470a",
  1967 => x"00000000",
  1968 => x"5374725f",
  1969 => x"325f4c6f",
  1970 => x"633a2020",
  1971 => x"20202020",
  1972 => x"20202020",
  1973 => x"2025730a",
  1974 => x"00000000",
  1975 => x"20202020",
  1976 => x"20202020",
  1977 => x"73686f75",
  1978 => x"6c642062",
  1979 => x"653a2020",
  1980 => x"20444852",
  1981 => x"5953544f",
  1982 => x"4e452050",
  1983 => x"524f4752",
  1984 => x"414d2c20",
  1985 => x"32274e44",
  1986 => x"20535452",
  1987 => x"494e470a",
  1988 => x"00000000",
  1989 => x"55736572",
  1990 => x"2074696d",
  1991 => x"653a2025",
  1992 => x"640a0000",
  1993 => x"4d696372",
  1994 => x"6f736563",
  1995 => x"6f6e6473",
  1996 => x"20666f72",
  1997 => x"206f6e65",
  1998 => x"2072756e",
  1999 => x"20746872",
  2000 => x"6f756768",
  2001 => x"20446872",
  2002 => x"7973746f",
  2003 => x"6e653a20",
  2004 => x"00000000",
  2005 => x"2564200a",
  2006 => x"00000000",
  2007 => x"44687279",
  2008 => x"73746f6e",
  2009 => x"65732070",
  2010 => x"65722053",
  2011 => x"65636f6e",
  2012 => x"643a2020",
  2013 => x"20202020",
  2014 => x"20202020",
  2015 => x"20202020",
  2016 => x"20202020",
  2017 => x"20202020",
  2018 => x"00000000",
  2019 => x"56415820",
  2020 => x"4d495053",
  2021 => x"20726174",
  2022 => x"696e6720",
  2023 => x"2a203130",
  2024 => x"3030203d",
  2025 => x"20256420",
  2026 => x"0a000000",
  2027 => x"50726f67",
  2028 => x"72616d20",
  2029 => x"636f6d70",
  2030 => x"696c6564",
  2031 => x"20776974",
  2032 => x"686f7574",
  2033 => x"20277265",
  2034 => x"67697374",
  2035 => x"65722720",
  2036 => x"61747472",
  2037 => x"69627574",
  2038 => x"650a0000",
  2039 => x"4d656173",
  2040 => x"75726564",
  2041 => x"2074696d",
  2042 => x"6520746f",
  2043 => x"6f20736d",
  2044 => x"616c6c20",
  2045 => x"746f206f",
  2046 => x"62746169",
  2047 => x"6e206d65",
  2048 => x"616e696e",
  2049 => x"6766756c",
  2050 => x"20726573",
  2051 => x"756c7473",
  2052 => x"0a000000",
  2053 => x"506c6561",
  2054 => x"73652069",
  2055 => x"6e637265",
  2056 => x"61736520",
  2057 => x"6e756d62",
  2058 => x"6572206f",
  2059 => x"66207275",
  2060 => x"6e730a00",
  2061 => x"44485259",
  2062 => x"53544f4e",
  2063 => x"45205052",
  2064 => x"4f475241",
  2065 => x"4d2c2033",
  2066 => x"27524420",
  2067 => x"53545249",
  2068 => x"4e470000",
  2069 => x"30313233",
  2070 => x"34353637",
  2071 => x"38394142",
  2072 => x"43444546",
  2073 => x"00000000",
  2074 => x"64756d6d",
  2075 => x"792e6578",
  2076 => x"65000000",
  2077 => x"43000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00002420",
  2082 => x"000061a8",
  2083 => x"00000000",
  2084 => x"00002068",
  2085 => x"00002098",
  2086 => x"00000000",
  2087 => x"00002300",
  2088 => x"0000235c",
  2089 => x"000023b8",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00002074",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000000",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000001",
  2129 => x"330eabcd",
  2130 => x"1234e66d",
  2131 => x"deec0005",
  2132 => x"000b0000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"00000000",
  2209 => x"00000000",
  2210 => x"00000000",
  2211 => x"00000000",
  2212 => x"00000000",
  2213 => x"00000000",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"00000000",
  2217 => x"00000000",
  2218 => x"00000000",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000000",
  2244 => x"00000000",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"00000000",
  2262 => x"00000000",
  2263 => x"00000000",
  2264 => x"00000000",
  2265 => x"00000000",
  2266 => x"00000000",
  2267 => x"00000000",
  2268 => x"00000000",
  2269 => x"00000000",
  2270 => x"00000000",
  2271 => x"00000000",
  2272 => x"00000000",
  2273 => x"00000000",
  2274 => x"00000000",
  2275 => x"00000000",
  2276 => x"00000000",
  2277 => x"00000000",
  2278 => x"00000000",
  2279 => x"00000000",
  2280 => x"00000000",
  2281 => x"00000000",
  2282 => x"00000000",
  2283 => x"00000000",
  2284 => x"00000000",
  2285 => x"00000000",
  2286 => x"00000000",
  2287 => x"00000000",
  2288 => x"00000000",
  2289 => x"00000000",
  2290 => x"00000000",
  2291 => x"00000000",
  2292 => x"00000000",
  2293 => x"00000000",
  2294 => x"00000000",
  2295 => x"00000000",
  2296 => x"00000000",
  2297 => x"00000000",
  2298 => x"00000000",
  2299 => x"00000000",
  2300 => x"00000000",
  2301 => x"00000000",
  2302 => x"00000000",
  2303 => x"00000000",
  2304 => x"00000000",
  2305 => x"00000000",
  2306 => x"00000000",
  2307 => x"00000000",
  2308 => x"00000000",
  2309 => x"ffffffff",
  2310 => x"00000000",
  2311 => x"ffffffff",
  2312 => x"00000000",
  2313 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;


-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b90",
     1 => x"fb040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"d3040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c9040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88ac",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba0",
   162 => x"ec738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88af0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b89",
   169 => x"9c040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"e5040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0ba1900c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"0b0b0b85",
   257 => x"8c3f0b0b",
   258 => x"0b98a83f",
   259 => x"04101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101010",
   266 => x"10101010",
   267 => x"53510473",
   268 => x"81ff0673",
   269 => x"83060981",
   270 => x"05830510",
   271 => x"10102b07",
   272 => x"72fc060c",
   273 => x"5151043c",
   274 => x"04727280",
   275 => x"728106ff",
   276 => x"05097206",
   277 => x"05711052",
   278 => x"720a100a",
   279 => x"5372ed38",
   280 => x"51515351",
   281 => x"040b0b0b",
   282 => x"0b80080b",
   283 => x"0b0b0b84",
   284 => x"080b0b0b",
   285 => x"0b880875",
   286 => x"750b0b0b",
   287 => x"8fa62d50",
   288 => x"500b0b0b",
   289 => x"0b800856",
   290 => x"0b0b0b0b",
   291 => x"880c0b0b",
   292 => x"0b0b840c",
   293 => x"0b0b0b0b",
   294 => x"800c5104",
   295 => x"0b0b0b0b",
   296 => x"80080b0b",
   297 => x"0b0b8408",
   298 => x"0b0b0b0b",
   299 => x"88087575",
   300 => x"0b0b0b8e",
   301 => x"bb2d5050",
   302 => x"0b0b0b0b",
   303 => x"8008560b",
   304 => x"0b0b0b88",
   305 => x"0c0b0b0b",
   306 => x"0b840c0b",
   307 => x"0b0b0b80",
   308 => x"0c51040b",
   309 => x"0b0b0b80",
   310 => x"080b0b0b",
   311 => x"0b84080b",
   312 => x"0b0b0b88",
   313 => x"080b0b0b",
   314 => x"91f42d0b",
   315 => x"0b0b0b88",
   316 => x"0c0b0b0b",
   317 => x"0b840c0b",
   318 => x"0b0b0b80",
   319 => x"0c04fe3d",
   320 => x"0d0b0b0b",
   321 => x"a8b80853",
   322 => x"84130870",
   323 => x"882a7081",
   324 => x"06515252",
   325 => x"70802e0b",
   326 => x"0b0b0bec",
   327 => x"387181ff",
   328 => x"060b0b0b",
   329 => x"0b800c84",
   330 => x"3d0d04ff",
   331 => x"3d0d0b0b",
   332 => x"0ba8b808",
   333 => x"52710870",
   334 => x"882a8132",
   335 => x"70810651",
   336 => x"5151700b",
   337 => x"0b0b0bed",
   338 => x"3873720c",
   339 => x"833d0d04",
   340 => x"0b0b0ba1",
   341 => x"9008802e",
   342 => x"0b0b0b0b",
   343 => x"ae380b0b",
   344 => x"0ba19408",
   345 => x"822e0b0b",
   346 => x"0b80c538",
   347 => x"8380800b",
   348 => x"0b0b0ba8",
   349 => x"b80c82a0",
   350 => x"800b0b0b",
   351 => x"0ba8bc0c",
   352 => x"8290800b",
   353 => x"0b0b0ba8",
   354 => x"c00c04f8",
   355 => x"808080a4",
   356 => x"0b0b0b0b",
   357 => x"a8b80cf8",
   358 => x"80808280",
   359 => x"0b0b0b0b",
   360 => x"a8bc0cf8",
   361 => x"80808480",
   362 => x"0b0b0b0b",
   363 => x"a8c00c04",
   364 => x"80c0a880",
   365 => x"8c0b0b0b",
   366 => x"0ba8b80c",
   367 => x"80c0a880",
   368 => x"940b0b0b",
   369 => x"0ba8bc0c",
   370 => x"0b0b0ba0",
   371 => x"fc0b0b0b",
   372 => x"0ba8c00c",
   373 => x"04f23d0d",
   374 => x"600b0b0b",
   375 => x"a8bc0856",
   376 => x"5d82750c",
   377 => x"8059805a",
   378 => x"800b8f3d",
   379 => x"5d5b7a10",
   380 => x"10157008",
   381 => x"7108719f",
   382 => x"2c7e852b",
   383 => x"5855557d",
   384 => x"5359570b",
   385 => x"0b0b81d9",
   386 => x"3f7d7f7a",
   387 => x"72077c72",
   388 => x"07717160",
   389 => x"8105415f",
   390 => x"5d5b5957",
   391 => x"55817b27",
   392 => x"0b0b0b0b",
   393 => x"9338767d",
   394 => x"0c77841e",
   395 => x"0c7c0b0b",
   396 => x"0b0b800c",
   397 => x"903d0d04",
   398 => x"0b0b0ba8",
   399 => x"bc08550b",
   400 => x"0b0bffaa",
   401 => x"39ff3d0d",
   402 => x"0b0b0ba8",
   403 => x"c4335170",
   404 => x"0b0b0b0b",
   405 => x"b7380b0b",
   406 => x"0ba19c08",
   407 => x"70085252",
   408 => x"70802e0b",
   409 => x"0b0b0b9c",
   410 => x"3884120b",
   411 => x"0b0ba19c",
   412 => x"0c702d0b",
   413 => x"0b0ba19c",
   414 => x"08700852",
   415 => x"52700b0b",
   416 => x"0b0be638",
   417 => x"810b0b0b",
   418 => x"0ba8c434",
   419 => x"833d0d04",
   420 => x"04803d0d",
   421 => x"0b0b0ba8",
   422 => x"b408802e",
   423 => x"0b0b0b0b",
   424 => x"92380b0b",
   425 => x"0b0b800b",
   426 => x"802e0981",
   427 => x"060b0b0b",
   428 => x"0b853882",
   429 => x"3d0d040b",
   430 => x"0b0ba8b4",
   431 => x"510b0b0b",
   432 => x"f2be3f82",
   433 => x"3d0d0404",
   434 => x"ff3d0d80",
   435 => x"52718113",
   436 => x"53ff800c",
   437 => x"71811353",
   438 => x"ff800c0b",
   439 => x"0b0b0bed",
   440 => x"39f93d0d",
   441 => x"797b7d7f",
   442 => x"56545254",
   443 => x"72802e0b",
   444 => x"0b0b0ba4",
   445 => x"38705771",
   446 => x"58a07331",
   447 => x"52807225",
   448 => x"0b0b0b0b",
   449 => x"a5387670",
   450 => x"742b5670",
   451 => x"732a7975",
   452 => x"2b075751",
   453 => x"74765351",
   454 => x"70740c71",
   455 => x"84150c73",
   456 => x"0b0b0b0b",
   457 => x"800c893d",
   458 => x"0d048055",
   459 => x"7672302b",
   460 => x"56747653",
   461 => x"510b0b0b",
   462 => x"0bde39fb",
   463 => x"3d0d7779",
   464 => x"55558056",
   465 => x"7575240b",
   466 => x"0b0b80c6",
   467 => x"38807424",
   468 => x"0b0b0b0b",
   469 => x"b0388053",
   470 => x"73527451",
   471 => x"0b0b0b81",
   472 => x"993f0b0b",
   473 => x"0b0b8008",
   474 => x"5475802e",
   475 => x"0b0b0b0b",
   476 => x"89380b0b",
   477 => x"0b0b8008",
   478 => x"3054730b",
   479 => x"0b0b0b80",
   480 => x"0c873d0d",
   481 => x"04733076",
   482 => x"81325754",
   483 => x"0b0b0b0b",
   484 => x"c5397430",
   485 => x"55815673",
   486 => x"80250b0b",
   487 => x"0bffb738",
   488 => x"0b0b0b0b",
   489 => x"e039fa3d",
   490 => x"0d787a57",
   491 => x"55805776",
   492 => x"75240b0b",
   493 => x"0b0bb838",
   494 => x"759f2c54",
   495 => x"81537574",
   496 => x"32743152",
   497 => x"74510b0b",
   498 => x"0b0baf3f",
   499 => x"0b0b0b0b",
   500 => x"80085476",
   501 => x"802e0b0b",
   502 => x"0b0b8938",
   503 => x"0b0b0b0b",
   504 => x"80083054",
   505 => x"730b0b0b",
   506 => x"0b800c88",
   507 => x"3d0d0474",
   508 => x"30558157",
   509 => x"0b0b0bff",
   510 => x"bf39fc3d",
   511 => x"0d767853",
   512 => x"54815380",
   513 => x"74732652",
   514 => x"5572802e",
   515 => x"0b0b0b0b",
   516 => x"a4387080",
   517 => x"2e0b0b0b",
   518 => x"0bb93880",
   519 => x"72240b0b",
   520 => x"0b0bb038",
   521 => x"71107310",
   522 => x"75722653",
   523 => x"5452720b",
   524 => x"0b0b0bde",
   525 => x"38735178",
   526 => x"0b0b0b0b",
   527 => x"83387451",
   528 => x"700b0b0b",
   529 => x"0b800c86",
   530 => x"3d0d0472",
   531 => x"812a7281",
   532 => x"2a535372",
   533 => x"802e0b0b",
   534 => x"0b0bda38",
   535 => x"7174260b",
   536 => x"0b0b0be7",
   537 => x"38737231",
   538 => x"75740774",
   539 => x"812a7481",
   540 => x"2a555556",
   541 => x"540b0b0b",
   542 => x"0bd939fd",
   543 => x"3d0d800b",
   544 => x"0b0b0ba1",
   545 => x"94085454",
   546 => x"72812e0b",
   547 => x"0b0b0baf",
   548 => x"38730b0b",
   549 => x"0ba8c80c",
   550 => x"0b0b0bf9",
   551 => x"b33f0b0b",
   552 => x"0bf6dd3f",
   553 => x"0b0b0ba1",
   554 => x"a0528151",
   555 => x"0b0b0bfc",
   556 => x"973f0b0b",
   557 => x"0b0b8008",
   558 => x"510b0b0b",
   559 => x"8af73f72",
   560 => x"0b0b0ba8",
   561 => x"c80c0b0b",
   562 => x"0bf9853f",
   563 => x"0b0b0bf6",
   564 => x"af3f0b0b",
   565 => x"0ba1a052",
   566 => x"81510b0b",
   567 => x"0bfbe93f",
   568 => x"0b0b0b0b",
   569 => x"8008510b",
   570 => x"0b0b8ac9",
   571 => x"3f000b0b",
   572 => x"0b0bfb39",
   573 => x"000b0b0b",
   574 => x"0bfb39f5",
   575 => x"3d0d7e60",
   576 => x"0b0b0ba8",
   577 => x"c808705b",
   578 => x"585b5b75",
   579 => x"0b0b0b80",
   580 => x"df38777a",
   581 => x"250b0b0b",
   582 => x"0bac3877",
   583 => x"1b703370",
   584 => x"81ff0658",
   585 => x"5859758a",
   586 => x"2e0b0b0b",
   587 => x"0ba33876",
   588 => x"81ff0651",
   589 => x"0b0b0bf7",
   590 => x"f23f8118",
   591 => x"58797824",
   592 => x"0b0b0b0b",
   593 => x"d638790b",
   594 => x"0b0b0b80",
   595 => x"0c8d3d0d",
   596 => x"048d510b",
   597 => x"0b0bf7d3",
   598 => x"3f783370",
   599 => x"81ff0652",
   600 => x"570b0b0b",
   601 => x"f7c53f81",
   602 => x"18580b0b",
   603 => x"0b0bce39",
   604 => x"79557a54",
   605 => x"7d538552",
   606 => x"8d3dfc05",
   607 => x"510b0b0b",
   608 => x"f5c53f0b",
   609 => x"0b0b0b80",
   610 => x"08560b0b",
   611 => x"0b89993f",
   612 => x"7b0b0b0b",
   613 => x"0b80080c",
   614 => x"750b0b0b",
   615 => x"0b800c8d",
   616 => x"3d0d04f6",
   617 => x"3d0d7d7f",
   618 => x"0b0b0ba8",
   619 => x"c808705b",
   620 => x"585a5a75",
   621 => x"0b0b0b80",
   622 => x"de387779",
   623 => x"250b0b0b",
   624 => x"80c8380b",
   625 => x"0b0bf6b6",
   626 => x"3f0b0b0b",
   627 => x"0b800881",
   628 => x"ff06708d",
   629 => x"32703070",
   630 => x"9f2a5151",
   631 => x"5757768a",
   632 => x"2e0b0b0b",
   633 => x"80e43875",
   634 => x"802e0b0b",
   635 => x"0b80db38",
   636 => x"771a5676",
   637 => x"76347651",
   638 => x"0b0b0bf6",
   639 => x"ae3f8118",
   640 => x"58787824",
   641 => x"0b0b0bff",
   642 => x"ba387756",
   643 => x"750b0b0b",
   644 => x"0b800c8c",
   645 => x"3d0d0478",
   646 => x"5579547c",
   647 => x"5384528c",
   648 => x"3dfc0551",
   649 => x"0b0b0bf4",
   650 => x"9e3f0b0b",
   651 => x"0b0b8008",
   652 => x"560b0b0b",
   653 => x"87f23f7a",
   654 => x"0b0b0b0b",
   655 => x"80080c75",
   656 => x"0b0b0b0b",
   657 => x"800c8c3d",
   658 => x"0d04771a",
   659 => x"568a7634",
   660 => x"8118588d",
   661 => x"510b0b0b",
   662 => x"f5d13f8a",
   663 => x"510b0b0b",
   664 => x"f5c93f77",
   665 => x"560b0b0b",
   666 => x"ffa239f9",
   667 => x"3d0d7957",
   668 => x"0b0b0ba8",
   669 => x"c808802e",
   670 => x"0b0b0b80",
   671 => x"c5387651",
   672 => x"0b0b0b8a",
   673 => x"b73f7b56",
   674 => x"7a550b0b",
   675 => x"0b0b8008",
   676 => x"81055476",
   677 => x"53825289",
   678 => x"3dfc0551",
   679 => x"0b0b0bf3",
   680 => x"a63f0b0b",
   681 => x"0b0b8008",
   682 => x"570b0b0b",
   683 => x"86fa3f77",
   684 => x"0b0b0b0b",
   685 => x"80080c76",
   686 => x"0b0b0b0b",
   687 => x"800c893d",
   688 => x"0d040b0b",
   689 => x"0b86e13f",
   690 => x"850b0b0b",
   691 => x"0b0b8008",
   692 => x"0cff0b0b",
   693 => x"0b0b0b80",
   694 => x"0c893d0d",
   695 => x"04fb3d0d",
   696 => x"0b0b0ba8",
   697 => x"c8087056",
   698 => x"54730b0b",
   699 => x"0b0b8c38",
   700 => x"740b0b0b",
   701 => x"0b800c87",
   702 => x"3d0d0477",
   703 => x"53835287",
   704 => x"3dfc0551",
   705 => x"0b0b0bf2",
   706 => x"be3f0b0b",
   707 => x"0b0b8008",
   708 => x"540b0b0b",
   709 => x"86923f75",
   710 => x"0b0b0b0b",
   711 => x"80080c73",
   712 => x"0b0b0b0b",
   713 => x"800c873d",
   714 => x"0d04ff0b",
   715 => x"0b0b0b0b",
   716 => x"800c04fb",
   717 => x"3d0d7755",
   718 => x"0b0b0ba8",
   719 => x"c808802e",
   720 => x"0b0b0b80",
   721 => x"c1387451",
   722 => x"0b0b0b88",
   723 => x"ef3f0b0b",
   724 => x"0b0b8008",
   725 => x"81055474",
   726 => x"53875287",
   727 => x"3dfc0551",
   728 => x"0b0b0bf1",
   729 => x"e23f0b0b",
   730 => x"0b0b8008",
   731 => x"550b0b0b",
   732 => x"85b63f75",
   733 => x"0b0b0b0b",
   734 => x"80080c74",
   735 => x"0b0b0b0b",
   736 => x"800c873d",
   737 => x"0d040b0b",
   738 => x"0b859d3f",
   739 => x"850b0b0b",
   740 => x"0b0b8008",
   741 => x"0cff0b0b",
   742 => x"0b0b0b80",
   743 => x"0c873d0d",
   744 => x"04fa3d0d",
   745 => x"0b0b0ba8",
   746 => x"c808802e",
   747 => x"0b0b0b0b",
   748 => x"b4387a55",
   749 => x"79547853",
   750 => x"8652883d",
   751 => x"fc05510b",
   752 => x"0b0bf183",
   753 => x"3f0b0b0b",
   754 => x"0b800856",
   755 => x"0b0b0b84",
   756 => x"d73f760b",
   757 => x"0b0b0b80",
   758 => x"080c750b",
   759 => x"0b0b0b80",
   760 => x"0c883d0d",
   761 => x"040b0b0b",
   762 => x"84be3f9d",
   763 => x"0b0b0b0b",
   764 => x"0b80080c",
   765 => x"ff0b0b0b",
   766 => x"0b0b800c",
   767 => x"883d0d04",
   768 => x"fb3d0d77",
   769 => x"79565680",
   770 => x"70545473",
   771 => x"75250b0b",
   772 => x"0b0ba338",
   773 => x"74101010",
   774 => x"f8055272",
   775 => x"16703370",
   776 => x"742b7607",
   777 => x"8116f816",
   778 => x"56565651",
   779 => x"51747324",
   780 => x"0b0b0b0b",
   781 => x"e638730b",
   782 => x"0b0b0b80",
   783 => x"0c873d0d",
   784 => x"04fc3d0d",
   785 => x"76785555",
   786 => x"bc538052",
   787 => x"73510b0b",
   788 => x"0b85b33f",
   789 => x"84527451",
   790 => x"0b0b0bff",
   791 => x"a33f0b0b",
   792 => x"0b0b8008",
   793 => x"74238452",
   794 => x"8415510b",
   795 => x"0b0bff90",
   796 => x"3f0b0b0b",
   797 => x"0b800882",
   798 => x"15238452",
   799 => x"8815510b",
   800 => x"0b0bfefc",
   801 => x"3f0b0b0b",
   802 => x"0b800884",
   803 => x"150c8452",
   804 => x"8c15510b",
   805 => x"0b0bfee8",
   806 => x"3f0b0b0b",
   807 => x"0b800888",
   808 => x"15238452",
   809 => x"9015510b",
   810 => x"0b0bfed4",
   811 => x"3f0b0b0b",
   812 => x"0b80088a",
   813 => x"15238452",
   814 => x"9415510b",
   815 => x"0b0bfec0",
   816 => x"3f0b0b0b",
   817 => x"0b80088c",
   818 => x"15238452",
   819 => x"9815510b",
   820 => x"0b0bfeac",
   821 => x"3f0b0b0b",
   822 => x"0b80088e",
   823 => x"15238852",
   824 => x"9c15510b",
   825 => x"0b0bfe98",
   826 => x"3f0b0b0b",
   827 => x"0b800890",
   828 => x"150c863d",
   829 => x"0d04e93d",
   830 => x"0d6a0b0b",
   831 => x"0ba8c808",
   832 => x"5757750b",
   833 => x"0b0b0b97",
   834 => x"3880c080",
   835 => x"0b84180c",
   836 => x"75ac180c",
   837 => x"750b0b0b",
   838 => x"0b800c99",
   839 => x"3d0d0489",
   840 => x"3d70556a",
   841 => x"54558a52",
   842 => x"993dffbc",
   843 => x"05510b0b",
   844 => x"0bee943f",
   845 => x"0b0b0b0b",
   846 => x"80087753",
   847 => x"7552560b",
   848 => x"0b0bfdfd",
   849 => x"3f0b0b0b",
   850 => x"81de3f77",
   851 => x"0b0b0b0b",
   852 => x"80080c75",
   853 => x"0b0b0b0b",
   854 => x"800c993d",
   855 => x"0d04e93d",
   856 => x"0d69570b",
   857 => x"0b0ba8c8",
   858 => x"08802e0b",
   859 => x"0b0b80d1",
   860 => x"3876510b",
   861 => x"0b0b84c4",
   862 => x"3f893d70",
   863 => x"560b0b0b",
   864 => x"0b800881",
   865 => x"05557754",
   866 => x"568f5299",
   867 => x"3dffbc05",
   868 => x"510b0b0b",
   869 => x"edb13f0b",
   870 => x"0b0b0b80",
   871 => x"086b5376",
   872 => x"52570b0b",
   873 => x"0bfd9a3f",
   874 => x"0b0b0b80",
   875 => x"fb3f770b",
   876 => x"0b0b0b80",
   877 => x"080c760b",
   878 => x"0b0b0b80",
   879 => x"0c993d0d",
   880 => x"040b0b0b",
   881 => x"80e23f85",
   882 => x"0b0b0b0b",
   883 => x"0b80080c",
   884 => x"ff0b0b0b",
   885 => x"0b0b800c",
   886 => x"993d0d04",
   887 => x"fc3d0d81",
   888 => x"540b0b0b",
   889 => x"a8c8080b",
   890 => x"0b0b0b8c",
   891 => x"38730b0b",
   892 => x"0b0b800c",
   893 => x"863d0d04",
   894 => x"765397b9",
   895 => x"52863dfc",
   896 => x"05510b0b",
   897 => x"0becc03f",
   898 => x"0b0b0b0b",
   899 => x"8008540b",
   900 => x"0b0b0b94",
   901 => x"3f740b0b",
   902 => x"0b0b8008",
   903 => x"0c730b0b",
   904 => x"0b0b800c",
   905 => x"863d0d04",
   906 => x"0b0b0ba1",
   907 => x"a4080b0b",
   908 => x"0b0b800c",
   909 => x"04f73d0d",
   910 => x"7b0b0b0b",
   911 => x"a1a40882",
   912 => x"c811085a",
   913 => x"545a7780",
   914 => x"2e0b0b0b",
   915 => x"80ee3881",
   916 => x"88188419",
   917 => x"08ff0581",
   918 => x"712b5955",
   919 => x"59807424",
   920 => x"0b0b0b81",
   921 => x"89388074",
   922 => x"240b0b0b",
   923 => x"0bbd3873",
   924 => x"822b7811",
   925 => x"88055656",
   926 => x"81801908",
   927 => x"77065372",
   928 => x"802e0b0b",
   929 => x"0b80c638",
   930 => x"78167008",
   931 => x"53537951",
   932 => x"74085372",
   933 => x"2dff14fc",
   934 => x"17fc1779",
   935 => x"812c5a57",
   936 => x"57547380",
   937 => x"250b0b0b",
   938 => x"0bce3877",
   939 => x"0858770b",
   940 => x"0b0bff9b",
   941 => x"380b0b0b",
   942 => x"a1a40853",
   943 => x"bc13080b",
   944 => x"0b0b0bb2",
   945 => x"3879510b",
   946 => x"0b0bf4a1",
   947 => x"3f740853",
   948 => x"722dff14",
   949 => x"fc17fc17",
   950 => x"79812c5a",
   951 => x"57575473",
   952 => x"80250b0b",
   953 => x"0bff9138",
   954 => x"0b0b0bff",
   955 => x"be398057",
   956 => x"0b0b0bfe",
   957 => x"f1397251",
   958 => x"bc130853",
   959 => x"722d7951",
   960 => x"0b0b0bf3",
   961 => x"e83ffc3d",
   962 => x"0d767971",
   963 => x"028c059f",
   964 => x"05335755",
   965 => x"53558372",
   966 => x"270b0b0b",
   967 => x"0b8e3874",
   968 => x"83065170",
   969 => x"802e0b0b",
   970 => x"0b0bae38",
   971 => x"ff125271",
   972 => x"ff2e0b0b",
   973 => x"0b0b9738",
   974 => x"73737081",
   975 => x"055534ff",
   976 => x"125271ff",
   977 => x"2e098106",
   978 => x"0b0b0b0b",
   979 => x"eb38740b",
   980 => x"0b0b0b80",
   981 => x"0c863d0d",
   982 => x"04747488",
   983 => x"2b750770",
   984 => x"71902b07",
   985 => x"5154518f",
   986 => x"72270b0b",
   987 => x"0b0ba938",
   988 => x"72717084",
   989 => x"05530c72",
   990 => x"71708405",
   991 => x"530c7271",
   992 => x"70840553",
   993 => x"0c727170",
   994 => x"8405530c",
   995 => x"f0125271",
   996 => x"8f260b0b",
   997 => x"0b0bd938",
   998 => x"8372270b",
   999 => x"0b0b0b94",
  1000 => x"38727170",
  1001 => x"8405530c",
  1002 => x"fc125271",
  1003 => x"83260b0b",
  1004 => x"0b0bee38",
  1005 => x"70530b0b",
  1006 => x"0bfef139",
  1007 => x"fd3d0d75",
  1008 => x"70718306",
  1009 => x"53555270",
  1010 => x"0b0b0b80",
  1011 => x"c0387170",
  1012 => x"087009f7",
  1013 => x"fbfdff12",
  1014 => x"0670f884",
  1015 => x"82818006",
  1016 => x"51515253",
  1017 => x"700b0b0b",
  1018 => x"0ba13884",
  1019 => x"13700870",
  1020 => x"09f7fbfd",
  1021 => x"ff120670",
  1022 => x"f8848281",
  1023 => x"80065151",
  1024 => x"52537080",
  1025 => x"2e0b0b0b",
  1026 => x"0be13872",
  1027 => x"52713351",
  1028 => x"70802e0b",
  1029 => x"0b0b0b8e",
  1030 => x"38811270",
  1031 => x"33525270",
  1032 => x"0b0b0b0b",
  1033 => x"f4387174",
  1034 => x"310b0b0b",
  1035 => x"0b800c85",
  1036 => x"3d0d04ff",
  1037 => x"3d0d0b0b",
  1038 => x"0ba8a80b",
  1039 => x"fc057008",
  1040 => x"525270ff",
  1041 => x"2e0b0b0b",
  1042 => x"0b953870",
  1043 => x"2dfc1270",
  1044 => x"08525270",
  1045 => x"ff2e0981",
  1046 => x"060b0b0b",
  1047 => x"0bed3883",
  1048 => x"3d0d0404",
  1049 => x"0b0b0beb",
  1050 => x"dc3f0400",
  1051 => x"00ffffff",
  1052 => x"ff00ffff",
  1053 => x"ffff00ff",
  1054 => x"ffffff00",
  1055 => x"00000040",
  1056 => x"64756d6d",
  1057 => x"792e6578",
  1058 => x"65000000",
  1059 => x"43000000",
  1060 => x"00000000",
  1061 => x"00000000",
  1062 => x"00000000",
  1063 => x"00001430",
  1064 => x"00001080",
  1065 => x"000010a8",
  1066 => x"00000000",
  1067 => x"00001310",
  1068 => x"0000136c",
  1069 => x"000013c8",
  1070 => x"00000000",
  1071 => x"00000000",
  1072 => x"00000000",
  1073 => x"00000000",
  1074 => x"00000000",
  1075 => x"00000000",
  1076 => x"00000000",
  1077 => x"00000000",
  1078 => x"00000000",
  1079 => x"0000108c",
  1080 => x"00000000",
  1081 => x"00000000",
  1082 => x"00000000",
  1083 => x"00000000",
  1084 => x"00000000",
  1085 => x"00000000",
  1086 => x"00000000",
  1087 => x"00000000",
  1088 => x"00000000",
  1089 => x"00000000",
  1090 => x"00000000",
  1091 => x"00000000",
  1092 => x"00000000",
  1093 => x"00000000",
  1094 => x"00000000",
  1095 => x"00000000",
  1096 => x"00000000",
  1097 => x"00000000",
  1098 => x"00000000",
  1099 => x"00000000",
  1100 => x"00000000",
  1101 => x"00000000",
  1102 => x"00000000",
  1103 => x"00000000",
  1104 => x"00000000",
  1105 => x"00000000",
  1106 => x"00000000",
  1107 => x"00000000",
  1108 => x"00000001",
  1109 => x"330eabcd",
  1110 => x"1234e66d",
  1111 => x"deec0005",
  1112 => x"000b0000",
  1113 => x"00000000",
  1114 => x"00000000",
  1115 => x"00000000",
  1116 => x"00000000",
  1117 => x"00000000",
  1118 => x"00000000",
  1119 => x"00000000",
  1120 => x"00000000",
  1121 => x"00000000",
  1122 => x"00000000",
  1123 => x"00000000",
  1124 => x"00000000",
  1125 => x"00000000",
  1126 => x"00000000",
  1127 => x"00000000",
  1128 => x"00000000",
  1129 => x"00000000",
  1130 => x"00000000",
  1131 => x"00000000",
  1132 => x"00000000",
  1133 => x"00000000",
  1134 => x"00000000",
  1135 => x"00000000",
  1136 => x"00000000",
  1137 => x"00000000",
  1138 => x"00000000",
  1139 => x"00000000",
  1140 => x"00000000",
  1141 => x"00000000",
  1142 => x"00000000",
  1143 => x"00000000",
  1144 => x"00000000",
  1145 => x"00000000",
  1146 => x"00000000",
  1147 => x"00000000",
  1148 => x"00000000",
  1149 => x"00000000",
  1150 => x"00000000",
  1151 => x"00000000",
  1152 => x"00000000",
  1153 => x"00000000",
  1154 => x"00000000",
  1155 => x"00000000",
  1156 => x"00000000",
  1157 => x"00000000",
  1158 => x"00000000",
  1159 => x"00000000",
  1160 => x"00000000",
  1161 => x"00000000",
  1162 => x"00000000",
  1163 => x"00000000",
  1164 => x"00000000",
  1165 => x"00000000",
  1166 => x"00000000",
  1167 => x"00000000",
  1168 => x"00000000",
  1169 => x"00000000",
  1170 => x"00000000",
  1171 => x"00000000",
  1172 => x"00000000",
  1173 => x"00000000",
  1174 => x"00000000",
  1175 => x"00000000",
  1176 => x"00000000",
  1177 => x"00000000",
  1178 => x"00000000",
  1179 => x"00000000",
  1180 => x"00000000",
  1181 => x"00000000",
  1182 => x"00000000",
  1183 => x"00000000",
  1184 => x"00000000",
  1185 => x"00000000",
  1186 => x"00000000",
  1187 => x"00000000",
  1188 => x"00000000",
  1189 => x"00000000",
  1190 => x"00000000",
  1191 => x"00000000",
  1192 => x"00000000",
  1193 => x"00000000",
  1194 => x"00000000",
  1195 => x"00000000",
  1196 => x"00000000",
  1197 => x"00000000",
  1198 => x"00000000",
  1199 => x"00000000",
  1200 => x"00000000",
  1201 => x"00000000",
  1202 => x"00000000",
  1203 => x"00000000",
  1204 => x"00000000",
  1205 => x"00000000",
  1206 => x"00000000",
  1207 => x"00000000",
  1208 => x"00000000",
  1209 => x"00000000",
  1210 => x"00000000",
  1211 => x"00000000",
  1212 => x"00000000",
  1213 => x"00000000",
  1214 => x"00000000",
  1215 => x"00000000",
  1216 => x"00000000",
  1217 => x"00000000",
  1218 => x"00000000",
  1219 => x"00000000",
  1220 => x"00000000",
  1221 => x"00000000",
  1222 => x"00000000",
  1223 => x"00000000",
  1224 => x"00000000",
  1225 => x"00000000",
  1226 => x"00000000",
  1227 => x"00000000",
  1228 => x"00000000",
  1229 => x"00000000",
  1230 => x"00000000",
  1231 => x"00000000",
  1232 => x"00000000",
  1233 => x"00000000",
  1234 => x"00000000",
  1235 => x"00000000",
  1236 => x"00000000",
  1237 => x"00000000",
  1238 => x"00000000",
  1239 => x"00000000",
  1240 => x"00000000",
  1241 => x"00000000",
  1242 => x"00000000",
  1243 => x"00000000",
  1244 => x"00000000",
  1245 => x"00000000",
  1246 => x"00000000",
  1247 => x"00000000",
  1248 => x"00000000",
  1249 => x"00000000",
  1250 => x"00000000",
  1251 => x"00000000",
  1252 => x"00000000",
  1253 => x"00000000",
  1254 => x"00000000",
  1255 => x"00000000",
  1256 => x"00000000",
  1257 => x"00000000",
  1258 => x"00000000",
  1259 => x"00000000",
  1260 => x"00000000",
  1261 => x"00000000",
  1262 => x"00000000",
  1263 => x"00000000",
  1264 => x"00000000",
  1265 => x"00000000",
  1266 => x"00000000",
  1267 => x"00000000",
  1268 => x"00000000",
  1269 => x"00000000",
  1270 => x"00000000",
  1271 => x"00000000",
  1272 => x"00000000",
  1273 => x"00000000",
  1274 => x"00000000",
  1275 => x"00000000",
  1276 => x"00000000",
  1277 => x"00000000",
  1278 => x"00000000",
  1279 => x"00000000",
  1280 => x"00000000",
  1281 => x"00000000",
  1282 => x"00000000",
  1283 => x"00000000",
  1284 => x"00000000",
  1285 => x"00000000",
  1286 => x"00000000",
  1287 => x"00000000",
  1288 => x"00000000",
  1289 => x"ffffffff",
  1290 => x"00000000",
  1291 => x"ffffffff",
  1292 => x"00000000",
  1293 => x"00000000",
  others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;

-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"f2040000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"95f87383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040ba0",
    29 => x"8080fd0b",
    30 => x"a08094f4",
    31 => x"040ba080",
    32 => x"80fd0402",
    33 => x"f8050d02",
    34 => x"8f05a080",
    35 => x"80b42d52",
    36 => x"ff840870",
    37 => x"882a7081",
    38 => x"06515151",
    39 => x"70802ef0",
    40 => x"3871ff84",
    41 => x"0c028805",
    42 => x"0d0402f4",
    43 => x"050d7453",
    44 => x"72a08080",
    45 => x"b42d7081",
    46 => x"ff065252",
    47 => x"70802ea3",
    48 => x"387181ff",
    49 => x"06811454",
    50 => x"52ff8408",
    51 => x"70882a70",
    52 => x"81065151",
    53 => x"5170802e",
    54 => x"f03871ff",
    55 => x"840ca080",
    56 => x"81b00402",
    57 => x"8c050d04",
    58 => x"02f8050d",
    59 => x"028f05a0",
    60 => x"8080b42d",
    61 => x"52ff8408",
    62 => x"70882a70",
    63 => x"81065151",
    64 => x"5170802e",
    65 => x"f03871ff",
    66 => x"840c0288",
    67 => x"050d0402",
    68 => x"d0050d02",
    69 => x"b405a080",
    70 => x"81e87170",
    71 => x"84055308",
    72 => x"5c5c5880",
    73 => x"7a708105",
    74 => x"5ca08080",
    75 => x"b42d5459",
    76 => x"72792e82",
    77 => x"cc3872a5",
    78 => x"2e098106",
    79 => x"82ab3879",
    80 => x"7081055b",
    81 => x"a08080b4",
    82 => x"2d537280",
    83 => x"e42e9f38",
    84 => x"7280e424",
    85 => x"8d387280",
    86 => x"e32e81c4",
    87 => x"38a08084",
    88 => x"b2047280",
    89 => x"f32e818d",
    90 => x"38a08084",
    91 => x"b2047784",
    92 => x"19710883",
    93 => x"ffe0e00b",
    94 => x"83ffe090",
    95 => x"595a5659",
    96 => x"53805673",
    97 => x"762e0981",
    98 => x"069538b0",
    99 => x"0b83ffe0",
   100 => x"900ba080",
   101 => x"80c92d81",
   102 => x"1555a080",
   103 => x"83c70473",
   104 => x"8f06a080",
   105 => x"96880553",
   106 => x"72a08080",
   107 => x"b42d7570",
   108 => x"810557a0",
   109 => x"8080c92d",
   110 => x"73842a54",
   111 => x"73e13874",
   112 => x"83ffe090",
   113 => x"2e9c38ff",
   114 => x"155574a0",
   115 => x"8080b42d",
   116 => x"77708105",
   117 => x"59a08080",
   118 => x"c92d8116",
   119 => x"56a08083",
   120 => x"bf048077",
   121 => x"a08080c9",
   122 => x"2d7583ff",
   123 => x"e0e05654",
   124 => x"a08084c6",
   125 => x"04778419",
   126 => x"71085759",
   127 => x"538075a0",
   128 => x"8080b42d",
   129 => x"54547274",
   130 => x"2ebc3881",
   131 => x"14701670",
   132 => x"a08080b4",
   133 => x"2d515454",
   134 => x"72f138a0",
   135 => x"8084c604",
   136 => x"77841983",
   137 => x"12a08080",
   138 => x"b42d5259",
   139 => x"53a08084",
   140 => x"e9048052",
   141 => x"a5517a2d",
   142 => x"80527251",
   143 => x"7a2d8219",
   144 => x"59a08084",
   145 => x"f20473ff",
   146 => x"15555380",
   147 => x"7325a338",
   148 => x"74708105",
   149 => x"56a08080",
   150 => x"b42d5380",
   151 => x"5272517a",
   152 => x"2d811959",
   153 => x"a08084c6",
   154 => x"04805272",
   155 => x"517a2d81",
   156 => x"19597970",
   157 => x"81055ba0",
   158 => x"8080b42d",
   159 => x"5372fdb6",
   160 => x"387883ff",
   161 => x"e0800c02",
   162 => x"b0050d04",
   163 => x"02f4050d",
   164 => x"74767181",
   165 => x"ff06c80c",
   166 => x"535383ff",
   167 => x"e1a00885",
   168 => x"3871892b",
   169 => x"5271982a",
   170 => x"c80c7190",
   171 => x"2a7081ff",
   172 => x"06c80c51",
   173 => x"71882a70",
   174 => x"81ff06c8",
   175 => x"0c517181",
   176 => x"ff06c80c",
   177 => x"72902a70",
   178 => x"81ff06c8",
   179 => x"0c51c808",
   180 => x"7081ff06",
   181 => x"515182b8",
   182 => x"bf527081",
   183 => x"ff2e0981",
   184 => x"06943881",
   185 => x"ff0bc80c",
   186 => x"c8087081",
   187 => x"ff06ff14",
   188 => x"54515171",
   189 => x"e5387083",
   190 => x"ffe0800c",
   191 => x"028c050d",
   192 => x"0402fc05",
   193 => x"0d81c751",
   194 => x"81ff0bc8",
   195 => x"0cff1151",
   196 => x"708025f4",
   197 => x"38028405",
   198 => x"0d0402f0",
   199 => x"050da080",
   200 => x"86812d81",
   201 => x"9c9f5380",
   202 => x"5287fc80",
   203 => x"f751a080",
   204 => x"858c2d83",
   205 => x"ffe08008",
   206 => x"5483ffe0",
   207 => x"8008812e",
   208 => x"098106ab",
   209 => x"3881ff0b",
   210 => x"c80c820a",
   211 => x"52849c80",
   212 => x"e951a080",
   213 => x"858c2d83",
   214 => x"ffe08008",
   215 => x"8d3881ff",
   216 => x"0bc80c73",
   217 => x"53a08086",
   218 => x"f604a080",
   219 => x"86812dff",
   220 => x"135372ff",
   221 => x"b2387283",
   222 => x"ffe0800c",
   223 => x"0290050d",
   224 => x"0402f405",
   225 => x"0d81ff0b",
   226 => x"c80c9353",
   227 => x"805287fc",
   228 => x"80c151a0",
   229 => x"80858c2d",
   230 => x"83ffe080",
   231 => x"088d3881",
   232 => x"ff0bc80c",
   233 => x"8153a080",
   234 => x"87b604a0",
   235 => x"8086812d",
   236 => x"ff135372",
   237 => x"d7387283",
   238 => x"ffe0800c",
   239 => x"028c050d",
   240 => x"0402f005",
   241 => x"0da08086",
   242 => x"812d83aa",
   243 => x"52849c80",
   244 => x"c851a080",
   245 => x"858c2d83",
   246 => x"ffe08008",
   247 => x"812e0981",
   248 => x"068e38cc",
   249 => x"0883ffff",
   250 => x"06537283",
   251 => x"aa2ea338",
   252 => x"a0808781",
   253 => x"2da08088",
   254 => x"8b048154",
   255 => x"a08089a2",
   256 => x"04a08096",
   257 => x"9c51a080",
   258 => x"828f2d80",
   259 => x"54a08089",
   260 => x"a20481ff",
   261 => x"0bc80cb1",
   262 => x"53a08086",
   263 => x"9a2d83ff",
   264 => x"e0800880",
   265 => x"2e80e238",
   266 => x"805287fc",
   267 => x"80fa51a0",
   268 => x"80858c2d",
   269 => x"83ffe080",
   270 => x"08bf3883",
   271 => x"ffe08008",
   272 => x"52a08096",
   273 => x"b851a080",
   274 => x"828f2d81",
   275 => x"ff0bc80c",
   276 => x"c80881ff",
   277 => x"067053a0",
   278 => x"8096c452",
   279 => x"54a08082",
   280 => x"8f2dcc08",
   281 => x"74862a70",
   282 => x"81067057",
   283 => x"51515372",
   284 => x"802eaf38",
   285 => x"a08087fa",
   286 => x"0483ffe0",
   287 => x"800852a0",
   288 => x"8096b851",
   289 => x"a080828f",
   290 => x"2d72822e",
   291 => x"fef338ff",
   292 => x"135372ff",
   293 => x"8438a080",
   294 => x"96d451a0",
   295 => x"8081aa2d",
   296 => x"72547383",
   297 => x"ffe0800c",
   298 => x"0290050d",
   299 => x"0402f405",
   300 => x"0d810b83",
   301 => x"ffe1a00c",
   302 => x"c408708f",
   303 => x"2a708106",
   304 => x"51515372",
   305 => x"f33872c4",
   306 => x"0ca08086",
   307 => x"812dc408",
   308 => x"708f2a70",
   309 => x"81065151",
   310 => x"5372f338",
   311 => x"810bc40c",
   312 => x"87538052",
   313 => x"84d480c0",
   314 => x"51a08085",
   315 => x"8c2d83ff",
   316 => x"e0800881",
   317 => x"2e098106",
   318 => x"873883ff",
   319 => x"e0800853",
   320 => x"a08096ec",
   321 => x"51a08081",
   322 => x"aa2d7282",
   323 => x"2e098106",
   324 => x"9238a080",
   325 => x"978051a0",
   326 => x"8081aa2d",
   327 => x"8053a080",
   328 => x"8b9304ff",
   329 => x"135372ff",
   330 => x"b938a080",
   331 => x"97a051a0",
   332 => x"8081aa2d",
   333 => x"a08087c1",
   334 => x"2d83ffe0",
   335 => x"800883ff",
   336 => x"e1a00c83",
   337 => x"ffe08008",
   338 => x"802e8b38",
   339 => x"a08097bc",
   340 => x"51a08081",
   341 => x"aa2da080",
   342 => x"97d051a0",
   343 => x"8081aa2d",
   344 => x"815287fc",
   345 => x"80d051a0",
   346 => x"80858c2d",
   347 => x"81ff0bc8",
   348 => x"0cc40870",
   349 => x"8f2a7081",
   350 => x"06515153",
   351 => x"72f33872",
   352 => x"c40c81ff",
   353 => x"0bc80ca0",
   354 => x"8097e051",
   355 => x"a08081aa",
   356 => x"2d815372",
   357 => x"83ffe080",
   358 => x"0c028c05",
   359 => x"0d04800b",
   360 => x"83ffe080",
   361 => x"0c0402e0",
   362 => x"050d797b",
   363 => x"57578058",
   364 => x"c408708f",
   365 => x"2a708106",
   366 => x"51515473",
   367 => x"f3388281",
   368 => x"0bc40c81",
   369 => x"ff0bc80c",
   370 => x"765287fc",
   371 => x"80d151a0",
   372 => x"80858c2d",
   373 => x"80dbc6df",
   374 => x"5583ffe0",
   375 => x"8008802e",
   376 => x"983883ff",
   377 => x"e0800853",
   378 => x"7652a080",
   379 => x"97ec51a0",
   380 => x"80828f2d",
   381 => x"a0808cc5",
   382 => x"0481ff0b",
   383 => x"c80cc808",
   384 => x"7081ff06",
   385 => x"51547381",
   386 => x"fe2e0981",
   387 => x"069b3880",
   388 => x"ff55cc08",
   389 => x"76708405",
   390 => x"580cff15",
   391 => x"55748025",
   392 => x"f1388158",
   393 => x"a0808caf",
   394 => x"04ff1555",
   395 => x"74cb3881",
   396 => x"ff0bc80c",
   397 => x"c408708f",
   398 => x"2a708106",
   399 => x"51515473",
   400 => x"f33873c4",
   401 => x"0c7783ff",
   402 => x"e0800c02",
   403 => x"a0050d04",
   404 => x"02f4050d",
   405 => x"7470882a",
   406 => x"83fe8006",
   407 => x"7072982a",
   408 => x"0772882b",
   409 => x"87fc8080",
   410 => x"0673982b",
   411 => x"81f00a06",
   412 => x"71730707",
   413 => x"83ffe080",
   414 => x"0c565153",
   415 => x"51028c05",
   416 => x"0d0402f4",
   417 => x"050d0292",
   418 => x"05227088",
   419 => x"2a71882b",
   420 => x"077083ff",
   421 => x"ff0683ff",
   422 => x"e0800c52",
   423 => x"52028c05",
   424 => x"0d0402f8",
   425 => x"050d7370",
   426 => x"902b7190",
   427 => x"2a0783ff",
   428 => x"e0800c52",
   429 => x"0288050d",
   430 => x"0402f405",
   431 => x"0d747652",
   432 => x"53807125",
   433 => x"90387052",
   434 => x"72708405",
   435 => x"5408ff13",
   436 => x"535171f4",
   437 => x"38028c05",
   438 => x"0d0402d8",
   439 => x"050d7b7d",
   440 => x"5b56810b",
   441 => x"a080988c",
   442 => x"59578359",
   443 => x"7708760c",
   444 => x"75087808",
   445 => x"56547375",
   446 => x"2e923875",
   447 => x"08537452",
   448 => x"a080989c",
   449 => x"51a08082",
   450 => x"8f2d8057",
   451 => x"79527551",
   452 => x"a0808db9",
   453 => x"2d750854",
   454 => x"73752e92",
   455 => x"38750853",
   456 => x"7452a080",
   457 => x"98dc51a0",
   458 => x"80828f2d",
   459 => x"8057ff19",
   460 => x"84195959",
   461 => x"788025ff",
   462 => x"b3387683",
   463 => x"ffe0800c",
   464 => x"02a8050d",
   465 => x"0402ec05",
   466 => x"0d765481",
   467 => x"5585aad5",
   468 => x"aad5740c",
   469 => x"fad5aad5",
   470 => x"aa0b8c15",
   471 => x"0ccc74a0",
   472 => x"8080c92d",
   473 => x"b30b8f15",
   474 => x"a08080c9",
   475 => x"2d730853",
   476 => x"72fce2d5",
   477 => x"aad52e90",
   478 => x"38730852",
   479 => x"a080999c",
   480 => x"51a08082",
   481 => x"8f2d8055",
   482 => x"8c140853",
   483 => x"72fad5aa",
   484 => x"d4b32e91",
   485 => x"388c1408",
   486 => x"52a08099",
   487 => x"d851a080",
   488 => x"828f2d80",
   489 => x"55775273",
   490 => x"51a0808d",
   491 => x"b92d7308",
   492 => x"5372fce2",
   493 => x"d5aad52e",
   494 => x"90387308",
   495 => x"52a0809a",
   496 => x"9451a080",
   497 => x"828f2d80",
   498 => x"558c1408",
   499 => x"5372fad5",
   500 => x"aad4b32e",
   501 => x"91388c14",
   502 => x"0852a080",
   503 => x"9ad051a0",
   504 => x"80828f2d",
   505 => x"80557483",
   506 => x"ffe0800c",
   507 => x"0294050d",
   508 => x"0402c805",
   509 => x"0d7f5c80",
   510 => x"0ba0809b",
   511 => x"8c525ba0",
   512 => x"80828f2d",
   513 => x"80e1b357",
   514 => x"8e5d7659",
   515 => x"8fffff5a",
   516 => x"76bfffff",
   517 => x"06771070",
   518 => x"962a7081",
   519 => x"06515758",
   520 => x"5874802e",
   521 => x"85387681",
   522 => x"07577695",
   523 => x"2a708106",
   524 => x"51557480",
   525 => x"2e853876",
   526 => x"81325776",
   527 => x"bfffff06",
   528 => x"7884291d",
   529 => x"79710c56",
   530 => x"7084291d",
   531 => x"56750c76",
   532 => x"1070962a",
   533 => x"70810651",
   534 => x"56577480",
   535 => x"2e853876",
   536 => x"81075776",
   537 => x"952a7081",
   538 => x"06515574",
   539 => x"802e8538",
   540 => x"76813257",
   541 => x"ff1a5a79",
   542 => x"8025ff94",
   543 => x"3878578f",
   544 => x"ffff5a76",
   545 => x"bfffff06",
   546 => x"77107096",
   547 => x"2a708106",
   548 => x"51575856",
   549 => x"74802e85",
   550 => x"38768107",
   551 => x"5776952a",
   552 => x"70810651",
   553 => x"5574802e",
   554 => x"85387681",
   555 => x"325776bf",
   556 => x"ffff0676",
   557 => x"84291d70",
   558 => x"08575a58",
   559 => x"74762ea7",
   560 => x"38807b53",
   561 => x"a0809ba0",
   562 => x"525ea080",
   563 => x"828f2d78",
   564 => x"08547553",
   565 => x"7552a080",
   566 => x"9bb451a0",
   567 => x"80828f2d",
   568 => x"7d5ba080",
   569 => x"91ea0481",
   570 => x"1b5b7784",
   571 => x"291c7008",
   572 => x"56567478",
   573 => x"2ea73880",
   574 => x"7b53a080",
   575 => x"9ba0525e",
   576 => x"a080828f",
   577 => x"2d750854",
   578 => x"77537752",
   579 => x"a0809bb4",
   580 => x"51a08082",
   581 => x"8f2d7d5b",
   582 => x"a08092a0",
   583 => x"04811b5b",
   584 => x"76107096",
   585 => x"2a708106",
   586 => x"51565774",
   587 => x"802e8538",
   588 => x"76810757",
   589 => x"76952a70",
   590 => x"81065155",
   591 => x"74802e85",
   592 => x"38768132",
   593 => x"57ff1a5a",
   594 => x"798025fe",
   595 => x"b638ff1d",
   596 => x"5d7cfdb6",
   597 => x"387d83ff",
   598 => x"e0800c02",
   599 => x"b8050d04",
   600 => x"02d0050d",
   601 => x"7d5b815a",
   602 => x"805980c0",
   603 => x"7a595c85",
   604 => x"ada989bb",
   605 => x"7b0c7957",
   606 => x"81569755",
   607 => x"77760782",
   608 => x"2b7b1151",
   609 => x"5485ada9",
   610 => x"89bb740c",
   611 => x"7510ff16",
   612 => x"56567480",
   613 => x"25e63877",
   614 => x"10811858",
   615 => x"58987725",
   616 => x"d7387e52",
   617 => x"7a51a080",
   618 => x"8db92d81",
   619 => x"58ff8787",
   620 => x"a5c37b0c",
   621 => x"97577782",
   622 => x"2b7b1170",
   623 => x"08565656",
   624 => x"73ff8787",
   625 => x"a5c32e09",
   626 => x"81068a38",
   627 => x"78780759",
   628 => x"a08093f2",
   629 => x"04740854",
   630 => x"7385ada9",
   631 => x"89bb2e92",
   632 => x"38807508",
   633 => x"547653a0",
   634 => x"809bdc52",
   635 => x"5aa08082",
   636 => x"8f2d7710",
   637 => x"ff185858",
   638 => x"768025ff",
   639 => x"b9387882",
   640 => x"2b597880",
   641 => x"2eb83878",
   642 => x"52a0809b",
   643 => x"fc51a080",
   644 => x"828f2d78",
   645 => x"992a8132",
   646 => x"70810670",
   647 => x"09810570",
   648 => x"72077009",
   649 => x"709f2c7f",
   650 => x"067e1087",
   651 => x"fffffe06",
   652 => x"62812c43",
   653 => x"5f5f5151",
   654 => x"56515578",
   655 => x"d6387909",
   656 => x"8105707b",
   657 => x"079f2a51",
   658 => x"547bbf24",
   659 => x"90387380",
   660 => x"2e8b38a0",
   661 => x"809c9451",
   662 => x"a080828f",
   663 => x"2d7b52a0",
   664 => x"809ce051",
   665 => x"a080828f",
   666 => x"2d7983ff",
   667 => x"e0800c02",
   668 => x"b0050d04",
   669 => x"02f8050d",
   670 => x"88bd0bff",
   671 => x"880ca080",
   672 => x"528051a0",
   673 => x"808dda2d",
   674 => x"83ffe080",
   675 => x"08802e8b",
   676 => x"38a0809d",
   677 => x"9c51a080",
   678 => x"828f2da0",
   679 => x"80528051",
   680 => x"a0808ec5",
   681 => x"2d83ffe0",
   682 => x"8008802e",
   683 => x"8b38a080",
   684 => x"9dc051a0",
   685 => x"80828f2d",
   686 => x"a0805280",
   687 => x"51a08092",
   688 => x"e02d83ff",
   689 => x"e0800880",
   690 => x"2e8b38a0",
   691 => x"809ddc51",
   692 => x"a080828f",
   693 => x"2d8051a0",
   694 => x"808ff12d",
   695 => x"83ffe080",
   696 => x"08802eff",
   697 => x"9938a080",
   698 => x"9df451a0",
   699 => x"80828f2d",
   700 => x"a08094fe",
   701 => x"04000000",
   702 => x"00ffffff",
   703 => x"ff00ffff",
   704 => x"ffff00ff",
   705 => x"ffffff00",
   706 => x"30313233",
   707 => x"34353637",
   708 => x"38394142",
   709 => x"43444546",
   710 => x"00000000",
   711 => x"53444843",
   712 => x"20496e69",
   713 => x"7469616c",
   714 => x"697a6174",
   715 => x"696f6e20",
   716 => x"6572726f",
   717 => x"72210a00",
   718 => x"434d4435",
   719 => x"38202564",
   720 => x"0a202000",
   721 => x"434d4435",
   722 => x"385f3220",
   723 => x"25640a20",
   724 => x"20000000",
   725 => x"44657465",
   726 => x"726d696e",
   727 => x"65642053",
   728 => x"44484320",
   729 => x"73746174",
   730 => x"75730a00",
   731 => x"53656e74",
   732 => x"20726573",
   733 => x"65742063",
   734 => x"6f6d6d61",
   735 => x"6e640a00",
   736 => x"53442063",
   737 => x"61726420",
   738 => x"696e6974",
   739 => x"69616c69",
   740 => x"7a617469",
   741 => x"6f6e2065",
   742 => x"72726f72",
   743 => x"210a0000",
   744 => x"43617264",
   745 => x"20726573",
   746 => x"706f6e64",
   747 => x"65642074",
   748 => x"6f207265",
   749 => x"7365740a",
   750 => x"00000000",
   751 => x"53444843",
   752 => x"20636172",
   753 => x"64206465",
   754 => x"74656374",
   755 => x"65640a00",
   756 => x"53656e64",
   757 => x"696e6720",
   758 => x"636d6431",
   759 => x"360a0000",
   760 => x"496e6974",
   761 => x"20646f6e",
   762 => x"650a0000",
   763 => x"52656164",
   764 => x"20636f6d",
   765 => x"6d616e64",
   766 => x"20666169",
   767 => x"6c656420",
   768 => x"61742025",
   769 => x"64202825",
   770 => x"64290a00",
   771 => x"00000000",
   772 => x"55555555",
   773 => x"aaaaaaaa",
   774 => x"ffffffff",
   775 => x"53616e69",
   776 => x"74792063",
   777 => x"6865636b",
   778 => x"20666169",
   779 => x"6c656420",
   780 => x"28626566",
   781 => x"6f726520",
   782 => x"63616368",
   783 => x"65207265",
   784 => x"66726573",
   785 => x"6829206f",
   786 => x"6e203078",
   787 => x"25642028",
   788 => x"676f7420",
   789 => x"30782564",
   790 => x"290a0000",
   791 => x"53616e69",
   792 => x"74792063",
   793 => x"6865636b",
   794 => x"20666169",
   795 => x"6c656420",
   796 => x"28616674",
   797 => x"65722063",
   798 => x"61636865",
   799 => x"20726566",
   800 => x"72657368",
   801 => x"29206f6e",
   802 => x"20307825",
   803 => x"64202867",
   804 => x"6f742030",
   805 => x"78256429",
   806 => x"0a000000",
   807 => x"42797465",
   808 => x"20636865",
   809 => x"636b2066",
   810 => x"61696c65",
   811 => x"64202862",
   812 => x"65666f72",
   813 => x"65206361",
   814 => x"63686520",
   815 => x"72656672",
   816 => x"65736829",
   817 => x"20617420",
   818 => x"30202867",
   819 => x"6f742030",
   820 => x"78256429",
   821 => x"0a000000",
   822 => x"42797465",
   823 => x"20636865",
   824 => x"636b2066",
   825 => x"61696c65",
   826 => x"64202862",
   827 => x"65666f72",
   828 => x"65206361",
   829 => x"63686520",
   830 => x"72656672",
   831 => x"65736829",
   832 => x"20617420",
   833 => x"33202867",
   834 => x"6f742030",
   835 => x"78256429",
   836 => x"0a000000",
   837 => x"42797465",
   838 => x"20636865",
   839 => x"636b2066",
   840 => x"61696c65",
   841 => x"64202861",
   842 => x"66746572",
   843 => x"20636163",
   844 => x"68652072",
   845 => x"65667265",
   846 => x"73682920",
   847 => x"61742030",
   848 => x"2028676f",
   849 => x"74203078",
   850 => x"2564290a",
   851 => x"00000000",
   852 => x"42797465",
   853 => x"20636865",
   854 => x"636b2066",
   855 => x"61696c65",
   856 => x"64202861",
   857 => x"66746572",
   858 => x"20636163",
   859 => x"68652072",
   860 => x"65667265",
   861 => x"73682920",
   862 => x"61742033",
   863 => x"2028676f",
   864 => x"74203078",
   865 => x"2564290a",
   866 => x"00000000",
   867 => x"43686563",
   868 => x"6b696e67",
   869 => x"206d656d",
   870 => x"6f72792e",
   871 => x"2e2e0a00",
   872 => x"30782564",
   873 => x"20676f6f",
   874 => x"64207265",
   875 => x"6164732c",
   876 => x"20000000",
   877 => x"4572726f",
   878 => x"72206174",
   879 => x"20307825",
   880 => x"642c2065",
   881 => x"78706563",
   882 => x"74656420",
   883 => x"30782564",
   884 => x"2c20676f",
   885 => x"74203078",
   886 => x"25640a00",
   887 => x"42616420",
   888 => x"64617461",
   889 => x"20666f75",
   890 => x"6e642061",
   891 => x"74203078",
   892 => x"25642028",
   893 => x"30782564",
   894 => x"290a0000",
   895 => x"416c6961",
   896 => x"73657320",
   897 => x"666f756e",
   898 => x"64206174",
   899 => x"20307825",
   900 => x"640a0000",
   901 => x"28416c69",
   902 => x"61736573",
   903 => x"2070726f",
   904 => x"6261626c",
   905 => x"79207369",
   906 => x"6d706c79",
   907 => x"20696e64",
   908 => x"69636174",
   909 => x"65207468",
   910 => x"61742052",
   911 => x"414d0a69",
   912 => x"7320736d",
   913 => x"616c6c65",
   914 => x"72207468",
   915 => x"616e2036",
   916 => x"34206d65",
   917 => x"67616279",
   918 => x"74657329",
   919 => x"0a000000",
   920 => x"53445241",
   921 => x"4d207369",
   922 => x"7a652028",
   923 => x"61737375",
   924 => x"6d696e67",
   925 => x"206e6f20",
   926 => x"61646472",
   927 => x"65737320",
   928 => x"6661756c",
   929 => x"74732920",
   930 => x"69732030",
   931 => x"78256420",
   932 => x"6d656761",
   933 => x"62797465",
   934 => x"730a0000",
   935 => x"46697273",
   936 => x"74207374",
   937 => x"61676520",
   938 => x"73616e69",
   939 => x"74792063",
   940 => x"6865636b",
   941 => x"20706173",
   942 => x"7365642e",
   943 => x"0a000000",
   944 => x"42797465",
   945 => x"20286471",
   946 => x"6d292063",
   947 => x"6865636b",
   948 => x"20706173",
   949 => x"7365640a",
   950 => x"00000000",
   951 => x"41646472",
   952 => x"65737320",
   953 => x"63686563",
   954 => x"6b207061",
   955 => x"73736564",
   956 => x"2e0a0000",
   957 => x"4c465352",
   958 => x"20636865",
   959 => x"636b2070",
   960 => x"61737365",
   961 => x"642e0a00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;


-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_ROM;

architecture arch of Dhrystone_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"80700b0b",
     2 => x"0bbfbc0c",
     3 => x"3a0b0b0b",
     4 => x"a8a90400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"8f040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bb3",
   162 => x"a4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f7040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"df040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bbfb80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"83dc3faa",
   257 => x"f43f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104b0",
   280 => x"08b408b8",
   281 => x"087575a2",
   282 => x"cf2d5050",
   283 => x"b00856b8",
   284 => x"0cb40cb0",
   285 => x"0c5104b0",
   286 => x"08b408b8",
   287 => x"087575a1",
   288 => x"9d2d5050",
   289 => x"b00856b8",
   290 => x"0cb40cb0",
   291 => x"0c5104b0",
   292 => x"08b408b8",
   293 => x"08a8ed2d",
   294 => x"b80cb40c",
   295 => x"b00c04fe",
   296 => x"3d0d0b0b",
   297 => x"80c6e808",
   298 => x"53841308",
   299 => x"70882a70",
   300 => x"81065152",
   301 => x"5270802e",
   302 => x"f0387181",
   303 => x"ff06b00c",
   304 => x"843d0d04",
   305 => x"ff3d0d0b",
   306 => x"0b80c6e8",
   307 => x"08527108",
   308 => x"70882a81",
   309 => x"32708106",
   310 => x"51515170",
   311 => x"f1387372",
   312 => x"0c833d0d",
   313 => x"04bfb808",
   314 => x"802ea338",
   315 => x"bfbc0882",
   316 => x"2ebd3883",
   317 => x"80800b0b",
   318 => x"0b80c6e8",
   319 => x"0c82a080",
   320 => x"0b80c6ec",
   321 => x"0c829080",
   322 => x"0b80c6f0",
   323 => x"0c04f880",
   324 => x"8080a40b",
   325 => x"0b0b80c6",
   326 => x"e80cf880",
   327 => x"8082800b",
   328 => x"80c6ec0c",
   329 => x"f8808084",
   330 => x"800b80c6",
   331 => x"f00c0480",
   332 => x"c0a8808c",
   333 => x"0b0b0b80",
   334 => x"c6e80c80",
   335 => x"c0a88094",
   336 => x"0b80c6ec",
   337 => x"0cb3b40b",
   338 => x"80c6f00c",
   339 => x"04f23d0d",
   340 => x"6080c6ec",
   341 => x"08565d82",
   342 => x"750c8059",
   343 => x"805a800b",
   344 => x"8f3d5d5b",
   345 => x"7a101015",
   346 => x"70087108",
   347 => x"719f2c7e",
   348 => x"852b5855",
   349 => x"557d5359",
   350 => x"5794ac3f",
   351 => x"7d7f7a72",
   352 => x"077c7207",
   353 => x"71716081",
   354 => x"05415f5d",
   355 => x"5b595755",
   356 => x"817b278f",
   357 => x"38767d0c",
   358 => x"77841e0c",
   359 => x"7cb00c90",
   360 => x"3d0d0480",
   361 => x"c6ec0855",
   362 => x"ffba39ff",
   363 => x"3d0d80c6",
   364 => x"f4335170",
   365 => x"a438bfc4",
   366 => x"08700852",
   367 => x"5270802e",
   368 => x"92388412",
   369 => x"bfc40c70",
   370 => x"2dbfc408",
   371 => x"70085252",
   372 => x"70f03881",
   373 => x"0b80c6f4",
   374 => x"34833d0d",
   375 => x"0404803d",
   376 => x"0d0b0b80",
   377 => x"c6e40880",
   378 => x"2e8e380b",
   379 => x"0b0b0b80",
   380 => x"0b802e09",
   381 => x"81068538",
   382 => x"823d0d04",
   383 => x"0b0b80c6",
   384 => x"e4510b0b",
   385 => x"0bf3f93f",
   386 => x"823d0d04",
   387 => x"04c008b0",
   388 => x"0c04803d",
   389 => x"0d80c10b",
   390 => x"81979834",
   391 => x"800b8199",
   392 => x"b00c70b0",
   393 => x"0c823d0d",
   394 => x"04ff3d0d",
   395 => x"800b8197",
   396 => x"98335252",
   397 => x"7080c12e",
   398 => x"99387181",
   399 => x"99b00807",
   400 => x"8199b00c",
   401 => x"80c20b81",
   402 => x"979c3470",
   403 => x"b00c833d",
   404 => x"0d04810b",
   405 => x"8199b008",
   406 => x"078199b0",
   407 => x"0c80c20b",
   408 => x"81979c34",
   409 => x"70b00c83",
   410 => x"3d0d04fd",
   411 => x"3d0d7570",
   412 => x"088a0553",
   413 => x"53819798",
   414 => x"33517080",
   415 => x"c12e8b38",
   416 => x"73f33870",
   417 => x"b00c853d",
   418 => x"0d04ff12",
   419 => x"70819794",
   420 => x"0831740c",
   421 => x"b00c853d",
   422 => x"0d04fc3d",
   423 => x"0d8197c0",
   424 => x"08557480",
   425 => x"2e8c3876",
   426 => x"7508710c",
   427 => x"8197c008",
   428 => x"56548c15",
   429 => x"53819794",
   430 => x"08528a51",
   431 => x"8c9c3f73",
   432 => x"b00c863d",
   433 => x"0d04fb3d",
   434 => x"0d777008",
   435 => x"5656b053",
   436 => x"8197c008",
   437 => x"52745198",
   438 => x"a23f850b",
   439 => x"8c170c85",
   440 => x"0b8c160c",
   441 => x"7508750c",
   442 => x"8197c008",
   443 => x"5473802e",
   444 => x"8a387308",
   445 => x"750c8197",
   446 => x"c008548c",
   447 => x"14538197",
   448 => x"9408528a",
   449 => x"518bd33f",
   450 => x"841508ad",
   451 => x"38860b8c",
   452 => x"160c8815",
   453 => x"52881608",
   454 => x"518adf3f",
   455 => x"8197c008",
   456 => x"7008760c",
   457 => x"548c1570",
   458 => x"54548a52",
   459 => x"7308518b",
   460 => x"a93f73b0",
   461 => x"0c873d0d",
   462 => x"04750854",
   463 => x"b0537352",
   464 => x"755197b7",
   465 => x"3f73b00c",
   466 => x"873d0d04",
   467 => x"f33d0d88",
   468 => x"bd0bff88",
   469 => x"0c8196ac",
   470 => x"0b8196e0",
   471 => x"0c8196e4",
   472 => x"0b8197c0",
   473 => x"0c8196ac",
   474 => x"0b8196e4",
   475 => x"0c800b81",
   476 => x"96e40b84",
   477 => x"050c820b",
   478 => x"8196e40b",
   479 => x"88050ca8",
   480 => x"0b8196e4",
   481 => x"0b8c050c",
   482 => x"9f53b3b8",
   483 => x"528196f4",
   484 => x"5196e83f",
   485 => x"9f53b3d8",
   486 => x"52819990",
   487 => x"5196dc3f",
   488 => x"8a0b80d4",
   489 => x"f80cbdfc",
   490 => x"518ddb3f",
   491 => x"b3f8518d",
   492 => x"d53fbdfc",
   493 => x"518dcf3f",
   494 => x"bfcc0880",
   495 => x"2e87ce38",
   496 => x"b4a8518d",
   497 => x"c13fbdfc",
   498 => x"518dbb3f",
   499 => x"bfc80852",
   500 => x"b4d4518d",
   501 => x"b13fc008",
   502 => x"80c8980c",
   503 => x"8158800b",
   504 => x"bfc80825",
   505 => x"82cf388c",
   506 => x"3d5b80c1",
   507 => x"0b819798",
   508 => x"34810b81",
   509 => x"99b00c80",
   510 => x"c20b8197",
   511 => x"9c34825c",
   512 => x"835a9f53",
   513 => x"b5845281",
   514 => x"97a05195",
   515 => x"ee3f815d",
   516 => x"800b8197",
   517 => x"a0538199",
   518 => x"9052558a",
   519 => x"e13fb008",
   520 => x"752e0981",
   521 => x"06833881",
   522 => x"55748199",
   523 => x"b00c7b70",
   524 => x"57557483",
   525 => x"25a03874",
   526 => x"101015fd",
   527 => x"055e8f3d",
   528 => x"fc055383",
   529 => x"52755189",
   530 => x"913f811c",
   531 => x"705d7057",
   532 => x"55837524",
   533 => x"e2387d54",
   534 => x"745380c8",
   535 => x"9c528197",
   536 => x"c8518986",
   537 => x"3f8197c0",
   538 => x"08700857",
   539 => x"57b05376",
   540 => x"52755195",
   541 => x"863f850b",
   542 => x"8c180c85",
   543 => x"0b8c170c",
   544 => x"7608760c",
   545 => x"8197c008",
   546 => x"5574802e",
   547 => x"8a387408",
   548 => x"760c8197",
   549 => x"c008558c",
   550 => x"15538197",
   551 => x"9408528a",
   552 => x"5188b73f",
   553 => x"84160887",
   554 => x"8b38860b",
   555 => x"8c170c88",
   556 => x"16528817",
   557 => x"085187c2",
   558 => x"3f8197c0",
   559 => x"08700877",
   560 => x"0c558c16",
   561 => x"7054578a",
   562 => x"52760851",
   563 => x"888c3f80",
   564 => x"c10b8197",
   565 => x"9c335656",
   566 => x"757526a2",
   567 => x"3880c352",
   568 => x"755188f0",
   569 => x"3fb0087d",
   570 => x"2e869c38",
   571 => x"81167081",
   572 => x"ff068197",
   573 => x"9c335757",
   574 => x"57747627",
   575 => x"e038797c",
   576 => x"297e7072",
   577 => x"35705f72",
   578 => x"72317087",
   579 => x"29723153",
   580 => x"538a0581",
   581 => x"97983381",
   582 => x"9794085a",
   583 => x"5a525b55",
   584 => x"7680c12e",
   585 => x"86a63878",
   586 => x"f7388118",
   587 => x"58bfc808",
   588 => x"7825fdb6",
   589 => x"38c00881",
   590 => x"96dc0cb5",
   591 => x"a4518ac6",
   592 => x"3fbdfc51",
   593 => x"8ac03fb5",
   594 => x"b4518aba",
   595 => x"3fbdfc51",
   596 => x"8ab43f81",
   597 => x"97940852",
   598 => x"b5ec518a",
   599 => x"a93f8552",
   600 => x"b688518a",
   601 => x"a13f8199",
   602 => x"b00852b6",
   603 => x"a4518a96",
   604 => x"3f8152b6",
   605 => x"88518a8e",
   606 => x"3f819798",
   607 => x"3352b6c0",
   608 => x"518a833f",
   609 => x"80c152b6",
   610 => x"dc5189fa",
   611 => x"3f81979c",
   612 => x"3352b6f8",
   613 => x"5189ef3f",
   614 => x"80c252b6",
   615 => x"dc5189e6",
   616 => x"3f8197e8",
   617 => x"0852b794",
   618 => x"5189db3f",
   619 => x"8752b688",
   620 => x"5189d33f",
   621 => x"80d4f808",
   622 => x"52b7b051",
   623 => x"89c83fb7",
   624 => x"cc5189c2",
   625 => x"3fb7f851",
   626 => x"89bc3f81",
   627 => x"97c00870",
   628 => x"085357b8",
   629 => x"845189ae",
   630 => x"3fb8a051",
   631 => x"89a83f81",
   632 => x"97c00884",
   633 => x"1108535b",
   634 => x"b8d45189",
   635 => x"993f8052",
   636 => x"b6885189",
   637 => x"913f8197",
   638 => x"c0088811",
   639 => x"085358b8",
   640 => x"f0518982",
   641 => x"3f8252b6",
   642 => x"885188fa",
   643 => x"3f8197c0",
   644 => x"088c1108",
   645 => x"5359b98c",
   646 => x"5188eb3f",
   647 => x"9152b688",
   648 => x"5188e33f",
   649 => x"8197c008",
   650 => x"900552b9",
   651 => x"a85188d6",
   652 => x"3fb9c451",
   653 => x"88d03fb9",
   654 => x"fc5188ca",
   655 => x"3f8196e0",
   656 => x"08700853",
   657 => x"55b88451",
   658 => x"88bc3fba",
   659 => x"905188b6",
   660 => x"3f8196e0",
   661 => x"08841108",
   662 => x"5356b8d4",
   663 => x"5188a73f",
   664 => x"8052b688",
   665 => x"51889f3f",
   666 => x"8196e008",
   667 => x"88110853",
   668 => x"57b8f051",
   669 => x"88903f81",
   670 => x"52b68851",
   671 => x"88883f81",
   672 => x"96e0088c",
   673 => x"1108535b",
   674 => x"b98c5187",
   675 => x"f93f9252",
   676 => x"b6885187",
   677 => x"f13f8196",
   678 => x"e0089005",
   679 => x"52b9a851",
   680 => x"87e43fb9",
   681 => x"c45187de",
   682 => x"3f7b52ba",
   683 => x"d05187d6",
   684 => x"3f8552b6",
   685 => x"885187ce",
   686 => x"3f7952ba",
   687 => x"ec5187c6",
   688 => x"3f8d52b6",
   689 => x"885187be",
   690 => x"3f7d52bb",
   691 => x"885187b6",
   692 => x"3f8752b6",
   693 => x"885187ae",
   694 => x"3f7c52bb",
   695 => x"a45187a6",
   696 => x"3f8152b6",
   697 => x"8851879e",
   698 => x"3f819990",
   699 => x"52bbc051",
   700 => x"87943fbb",
   701 => x"dc51878e",
   702 => x"3f8197a0",
   703 => x"52bc9451",
   704 => x"87843fbc",
   705 => x"b05186fe",
   706 => x"3fbdfc51",
   707 => x"86f83f81",
   708 => x"96dc0880",
   709 => x"c8980831",
   710 => x"7080c894",
   711 => x"0c52bce8",
   712 => x"5186e33f",
   713 => x"80c89408",
   714 => x"5680f776",
   715 => x"2580e438",
   716 => x"bfc80870",
   717 => x"7787e829",
   718 => x"3580c88c",
   719 => x"0c767187",
   720 => x"e8293580",
   721 => x"c8900c76",
   722 => x"7184b929",
   723 => x"358197c4",
   724 => x"0c5abcf8",
   725 => x"5186af3f",
   726 => x"80c88c08",
   727 => x"52bda851",
   728 => x"86a43fbd",
   729 => x"b051869e",
   730 => x"3f80c890",
   731 => x"0852bda8",
   732 => x"5186933f",
   733 => x"8197c408",
   734 => x"52bde051",
   735 => x"86883fbd",
   736 => x"fc518682",
   737 => x"3f800bb0",
   738 => x"0c8f3d0d",
   739 => x"04be8051",
   740 => x"f8b139be",
   741 => x"b05185ee",
   742 => x"3fbee851",
   743 => x"85e83fbd",
   744 => x"fc5185e2",
   745 => x"3f80c894",
   746 => x"08bfc808",
   747 => x"707287e8",
   748 => x"293580c8",
   749 => x"8c0c7171",
   750 => x"87e82935",
   751 => x"80c8900c",
   752 => x"717184b9",
   753 => x"29358197",
   754 => x"c40c5b56",
   755 => x"bcf85185",
   756 => x"b53f80c8",
   757 => x"8c0852bd",
   758 => x"a85185aa",
   759 => x"3fbdb051",
   760 => x"85a43f80",
   761 => x"c8900852",
   762 => x"bda85185",
   763 => x"993f8197",
   764 => x"c40852bd",
   765 => x"e051858e",
   766 => x"3fbdfc51",
   767 => x"85883f80",
   768 => x"0bb00c8f",
   769 => x"3d0d048f",
   770 => x"3df80552",
   771 => x"805180ea",
   772 => x"3f9f53bf",
   773 => x"88528197",
   774 => x"a0518ddf",
   775 => x"3f777881",
   776 => x"97940c81",
   777 => x"177081ff",
   778 => x"0681979c",
   779 => x"33585858",
   780 => x"5af9c639",
   781 => x"760856b0",
   782 => x"53755276",
   783 => x"518dbc3f",
   784 => x"80c10b81",
   785 => x"979c3356",
   786 => x"56f98d39",
   787 => x"ff157077",
   788 => x"317c0c59",
   789 => x"800b8119",
   790 => x"5959bfc8",
   791 => x"087825f7",
   792 => x"8938f9d1",
   793 => x"39ff3d0d",
   794 => x"73823270",
   795 => x"30707207",
   796 => x"8025b00c",
   797 => x"5252833d",
   798 => x"0d04fe3d",
   799 => x"0d747671",
   800 => x"53545271",
   801 => x"822e8338",
   802 => x"83517181",
   803 => x"2e9a3881",
   804 => x"72269f38",
   805 => x"71822eb8",
   806 => x"3871842e",
   807 => x"a9387073",
   808 => x"0c70b00c",
   809 => x"843d0d04",
   810 => x"80e40b81",
   811 => x"97940825",
   812 => x"8b388073",
   813 => x"0c70b00c",
   814 => x"843d0d04",
   815 => x"83730c70",
   816 => x"b00c843d",
   817 => x"0d048273",
   818 => x"0c70b00c",
   819 => x"843d0d04",
   820 => x"81730c70",
   821 => x"b00c843d",
   822 => x"0d04803d",
   823 => x"0d747414",
   824 => x"8205710c",
   825 => x"b00c823d",
   826 => x"0d04f73d",
   827 => x"0d7b7d7f",
   828 => x"61851270",
   829 => x"822b7511",
   830 => x"70747170",
   831 => x"8405530c",
   832 => x"5a5a5d5b",
   833 => x"760c7980",
   834 => x"f8180c79",
   835 => x"86125257",
   836 => x"585a5a76",
   837 => x"76249938",
   838 => x"76b32982",
   839 => x"2b791151",
   840 => x"53767370",
   841 => x"8405550c",
   842 => x"81145475",
   843 => x"7425f238",
   844 => x"7681cc29",
   845 => x"19fc1108",
   846 => x"8105fc12",
   847 => x"0c7a1970",
   848 => x"089fa013",
   849 => x"0c585685",
   850 => x"0b819794",
   851 => x"0c75b00c",
   852 => x"8b3d0d04",
   853 => x"fe3d0d02",
   854 => x"93053351",
   855 => x"80028405",
   856 => x"97053354",
   857 => x"5270732e",
   858 => x"883871b0",
   859 => x"0c843d0d",
   860 => x"04708197",
   861 => x"9834810b",
   862 => x"b00c843d",
   863 => x"0d04f83d",
   864 => x"0d7a7c59",
   865 => x"56820b83",
   866 => x"19555574",
   867 => x"16703375",
   868 => x"335b5153",
   869 => x"72792e80",
   870 => x"c63880c1",
   871 => x"0b811681",
   872 => x"16565657",
   873 => x"827525e3",
   874 => x"38ffa917",
   875 => x"7081ff06",
   876 => x"55597382",
   877 => x"26833887",
   878 => x"55815376",
   879 => x"80d22e98",
   880 => x"38775275",
   881 => x"518bcd3f",
   882 => x"805372b0",
   883 => x"08258938",
   884 => x"87158197",
   885 => x"940c8153",
   886 => x"72b00c8a",
   887 => x"3d0d0472",
   888 => x"81979834",
   889 => x"827525ff",
   890 => x"a238ffbd",
   891 => x"39ff3d0d",
   892 => x"7352ff84",
   893 => x"0870882a",
   894 => x"70810651",
   895 => x"51517080",
   896 => x"2ef03871",
   897 => x"ff840c71",
   898 => x"b00c833d",
   899 => x"0d04fd3d",
   900 => x"0d755380",
   901 => x"73335254",
   902 => x"70742ea4",
   903 => x"38705281",
   904 => x"1353ff84",
   905 => x"0870882a",
   906 => x"70810651",
   907 => x"51517080",
   908 => x"2ef03871",
   909 => x"ff840c81",
   910 => x"14733353",
   911 => x"5471e038",
   912 => x"73b00c85",
   913 => x"3d0d04ff",
   914 => x"3d0dff84",
   915 => x"0870892a",
   916 => x"70810651",
   917 => x"52527080",
   918 => x"2ef03871",
   919 => x"81ff06b0",
   920 => x"0c833d0d",
   921 => x"04fe3d0d",
   922 => x"74c00853",
   923 => x"5372802e",
   924 => x"9138c008",
   925 => x"5170722e",
   926 => x"f93870ff",
   927 => x"14545272",
   928 => x"f138843d",
   929 => x"0d04f13d",
   930 => x"0d923d80",
   931 => x"c7c85c5c",
   932 => x"807c7084",
   933 => x"055e0871",
   934 => x"5f5f587d",
   935 => x"7084055f",
   936 => x"0857805a",
   937 => x"76982a77",
   938 => x"882b5855",
   939 => x"74802e81",
   940 => x"ef387c80",
   941 => x"2eb73880",
   942 => x"5d7480e4",
   943 => x"2e819838",
   944 => x"7480e426",
   945 => x"80d83874",
   946 => x"80e32eb7",
   947 => x"38a551fe",
   948 => x"9c3f7451",
   949 => x"fe973f82",
   950 => x"1858811a",
   951 => x"5a837a25",
   952 => x"c33874ff",
   953 => x"b6387eb0",
   954 => x"0c913d0d",
   955 => x"0474a52e",
   956 => x"09810697",
   957 => x"38810b81",
   958 => x"1b5b5d83",
   959 => x"7a25ffa4",
   960 => x"38e0397b",
   961 => x"841d7108",
   962 => x"575d5474",
   963 => x"51fdde3f",
   964 => x"8118811b",
   965 => x"5b58837a",
   966 => x"25ff8938",
   967 => x"c5397480",
   968 => x"f32e0981",
   969 => x"06ffa638",
   970 => x"7b841d71",
   971 => x"0870545d",
   972 => x"5d53fdda",
   973 => x"3f800bff",
   974 => x"11545280",
   975 => x"7225ff9a",
   976 => x"387a7081",
   977 => x"055c3370",
   978 => x"5255fda1",
   979 => x"3f811873",
   980 => x"ff155553",
   981 => x"58e5397b",
   982 => x"841d7108",
   983 => x"7f5c555d",
   984 => x"52875672",
   985 => x"9c2a7384",
   986 => x"2b545271",
   987 => x"802e8338",
   988 => x"8159b712",
   989 => x"54718924",
   990 => x"8438b012",
   991 => x"54789238",
   992 => x"ff165675",
   993 => x"8025dc38",
   994 => x"800bff11",
   995 => x"5452ffab",
   996 => x"397351fc",
   997 => x"d83fff16",
   998 => x"56758025",
   999 => x"c638e939",
  1000 => x"77b00c91",
  1001 => x"3d0d04bc",
  1002 => x"0802bc0c",
  1003 => x"f53d0dbc",
  1004 => x"08940508",
  1005 => x"9d38bc08",
  1006 => x"8c0508bc",
  1007 => x"08900508",
  1008 => x"bc088805",
  1009 => x"08585654",
  1010 => x"73760c74",
  1011 => x"84170c81",
  1012 => x"bf39800b",
  1013 => x"bc08f005",
  1014 => x"0c800bbc",
  1015 => x"08f4050c",
  1016 => x"bc088c05",
  1017 => x"08bc0890",
  1018 => x"05085654",
  1019 => x"73bc08f0",
  1020 => x"050c74bc",
  1021 => x"08f4050c",
  1022 => x"bc08f805",
  1023 => x"bc08f005",
  1024 => x"56568870",
  1025 => x"54755376",
  1026 => x"525485ef",
  1027 => x"3fa00bbc",
  1028 => x"08940508",
  1029 => x"31bc08ec",
  1030 => x"050cbc08",
  1031 => x"ec050880",
  1032 => x"249d3880",
  1033 => x"0bbc08f4",
  1034 => x"050cbc08",
  1035 => x"ec050830",
  1036 => x"bc08fc05",
  1037 => x"08712bbc",
  1038 => x"08f0050c",
  1039 => x"54b939bc",
  1040 => x"08fc0508",
  1041 => x"bc08ec05",
  1042 => x"082abc08",
  1043 => x"e8050cbc",
  1044 => x"08fc0508",
  1045 => x"bc089405",
  1046 => x"082bbc08",
  1047 => x"f4050cbc",
  1048 => x"08f80508",
  1049 => x"bc089405",
  1050 => x"082b70bc",
  1051 => x"08e80508",
  1052 => x"07bc08f0",
  1053 => x"050c54bc",
  1054 => x"08f00508",
  1055 => x"bc08f405",
  1056 => x"08bc0888",
  1057 => x"05085856",
  1058 => x"5473760c",
  1059 => x"7484170c",
  1060 => x"bc088805",
  1061 => x"08b00c8d",
  1062 => x"3d0dbc0c",
  1063 => x"04bc0802",
  1064 => x"bc0cf93d",
  1065 => x"0d800bbc",
  1066 => x"08fc050c",
  1067 => x"bc088805",
  1068 => x"088025ab",
  1069 => x"38bc0888",
  1070 => x"050830bc",
  1071 => x"0888050c",
  1072 => x"800bbc08",
  1073 => x"f4050cbc",
  1074 => x"08fc0508",
  1075 => x"8838810b",
  1076 => x"bc08f405",
  1077 => x"0cbc08f4",
  1078 => x"0508bc08",
  1079 => x"fc050cbc",
  1080 => x"088c0508",
  1081 => x"8025ab38",
  1082 => x"bc088c05",
  1083 => x"0830bc08",
  1084 => x"8c050c80",
  1085 => x"0bbc08f0",
  1086 => x"050cbc08",
  1087 => x"fc050888",
  1088 => x"38810bbc",
  1089 => x"08f0050c",
  1090 => x"bc08f005",
  1091 => x"08bc08fc",
  1092 => x"050c8053",
  1093 => x"bc088c05",
  1094 => x"0852bc08",
  1095 => x"88050851",
  1096 => x"81a73fb0",
  1097 => x"0870bc08",
  1098 => x"f8050c54",
  1099 => x"bc08fc05",
  1100 => x"08802e8c",
  1101 => x"38bc08f8",
  1102 => x"050830bc",
  1103 => x"08f8050c",
  1104 => x"bc08f805",
  1105 => x"0870b00c",
  1106 => x"54893d0d",
  1107 => x"bc0c04bc",
  1108 => x"0802bc0c",
  1109 => x"fb3d0d80",
  1110 => x"0bbc08fc",
  1111 => x"050cbc08",
  1112 => x"88050880",
  1113 => x"259338bc",
  1114 => x"08880508",
  1115 => x"30bc0888",
  1116 => x"050c810b",
  1117 => x"bc08fc05",
  1118 => x"0cbc088c",
  1119 => x"05088025",
  1120 => x"8c38bc08",
  1121 => x"8c050830",
  1122 => x"bc088c05",
  1123 => x"0c8153bc",
  1124 => x"088c0508",
  1125 => x"52bc0888",
  1126 => x"050851ad",
  1127 => x"3fb00870",
  1128 => x"bc08f805",
  1129 => x"0c54bc08",
  1130 => x"fc050880",
  1131 => x"2e8c38bc",
  1132 => x"08f80508",
  1133 => x"30bc08f8",
  1134 => x"050cbc08",
  1135 => x"f8050870",
  1136 => x"b00c5487",
  1137 => x"3d0dbc0c",
  1138 => x"04bc0802",
  1139 => x"bc0cfd3d",
  1140 => x"0d810bbc",
  1141 => x"08fc050c",
  1142 => x"800bbc08",
  1143 => x"f8050cbc",
  1144 => x"088c0508",
  1145 => x"bc088805",
  1146 => x"0827ac38",
  1147 => x"bc08fc05",
  1148 => x"08802ea3",
  1149 => x"38800bbc",
  1150 => x"088c0508",
  1151 => x"249938bc",
  1152 => x"088c0508",
  1153 => x"10bc088c",
  1154 => x"050cbc08",
  1155 => x"fc050810",
  1156 => x"bc08fc05",
  1157 => x"0cc939bc",
  1158 => x"08fc0508",
  1159 => x"802e80c9",
  1160 => x"38bc088c",
  1161 => x"0508bc08",
  1162 => x"88050826",
  1163 => x"a138bc08",
  1164 => x"880508bc",
  1165 => x"088c0508",
  1166 => x"31bc0888",
  1167 => x"050cbc08",
  1168 => x"f80508bc",
  1169 => x"08fc0508",
  1170 => x"07bc08f8",
  1171 => x"050cbc08",
  1172 => x"fc050881",
  1173 => x"2abc08fc",
  1174 => x"050cbc08",
  1175 => x"8c050881",
  1176 => x"2abc088c",
  1177 => x"050cffaf",
  1178 => x"39bc0890",
  1179 => x"0508802e",
  1180 => x"8f38bc08",
  1181 => x"88050870",
  1182 => x"bc08f405",
  1183 => x"0c518d39",
  1184 => x"bc08f805",
  1185 => x"0870bc08",
  1186 => x"f4050c51",
  1187 => x"bc08f405",
  1188 => x"08b00c85",
  1189 => x"3d0dbc0c",
  1190 => x"04bc0802",
  1191 => x"bc0cff3d",
  1192 => x"0d800bbc",
  1193 => x"08fc050c",
  1194 => x"bc088805",
  1195 => x"088106ff",
  1196 => x"11700970",
  1197 => x"bc088c05",
  1198 => x"0806bc08",
  1199 => x"fc050811",
  1200 => x"bc08fc05",
  1201 => x"0cbc0888",
  1202 => x"0508812a",
  1203 => x"bc088805",
  1204 => x"0cbc088c",
  1205 => x"050810bc",
  1206 => x"088c050c",
  1207 => x"51515151",
  1208 => x"bc088805",
  1209 => x"08802e84",
  1210 => x"38ffbd39",
  1211 => x"bc08fc05",
  1212 => x"0870b00c",
  1213 => x"51833d0d",
  1214 => x"bc0c04fc",
  1215 => x"3d0d7670",
  1216 => x"797b5555",
  1217 => x"55558f72",
  1218 => x"278c3872",
  1219 => x"75078306",
  1220 => x"5170802e",
  1221 => x"a738ff12",
  1222 => x"5271ff2e",
  1223 => x"98387270",
  1224 => x"81055433",
  1225 => x"74708105",
  1226 => x"5634ff12",
  1227 => x"5271ff2e",
  1228 => x"098106ea",
  1229 => x"3874b00c",
  1230 => x"863d0d04",
  1231 => x"74517270",
  1232 => x"84055408",
  1233 => x"71708405",
  1234 => x"530c7270",
  1235 => x"84055408",
  1236 => x"71708405",
  1237 => x"530c7270",
  1238 => x"84055408",
  1239 => x"71708405",
  1240 => x"530c7270",
  1241 => x"84055408",
  1242 => x"71708405",
  1243 => x"530cf012",
  1244 => x"52718f26",
  1245 => x"c9388372",
  1246 => x"27953872",
  1247 => x"70840554",
  1248 => x"08717084",
  1249 => x"05530cfc",
  1250 => x"12527183",
  1251 => x"26ed3870",
  1252 => x"54ff8339",
  1253 => x"fb3d0d77",
  1254 => x"79707207",
  1255 => x"83065354",
  1256 => x"52709338",
  1257 => x"71737308",
  1258 => x"54565471",
  1259 => x"73082e80",
  1260 => x"c4387375",
  1261 => x"54527133",
  1262 => x"7081ff06",
  1263 => x"52547080",
  1264 => x"2e9d3872",
  1265 => x"33557075",
  1266 => x"2e098106",
  1267 => x"95388112",
  1268 => x"81147133",
  1269 => x"7081ff06",
  1270 => x"54565452",
  1271 => x"70e53872",
  1272 => x"33557381",
  1273 => x"ff067581",
  1274 => x"ff067171",
  1275 => x"31b00c52",
  1276 => x"52873d0d",
  1277 => x"04710970",
  1278 => x"f7fbfdff",
  1279 => x"140670f8",
  1280 => x"84828180",
  1281 => x"06515151",
  1282 => x"70973884",
  1283 => x"14841671",
  1284 => x"08545654",
  1285 => x"7175082e",
  1286 => x"dc387375",
  1287 => x"5452ff96",
  1288 => x"39800bb0",
  1289 => x"0c873d0d",
  1290 => x"04fd3d0d",
  1291 => x"800bbfbc",
  1292 => x"08545472",
  1293 => x"812e9a38",
  1294 => x"7380c888",
  1295 => x"0ce1a63f",
  1296 => x"dfbe3fbf",
  1297 => x"d0528151",
  1298 => x"e6823fb0",
  1299 => x"08518799",
  1300 => x"3f7280c8",
  1301 => x"880ce18d",
  1302 => x"3fdfa53f",
  1303 => x"bfd05281",
  1304 => x"51e5e93f",
  1305 => x"b0085187",
  1306 => x"803f00ff",
  1307 => x"3900ff39",
  1308 => x"f53d0d7e",
  1309 => x"6080c888",
  1310 => x"08705b58",
  1311 => x"5b5b7580",
  1312 => x"c238777a",
  1313 => x"25a13877",
  1314 => x"1b703370",
  1315 => x"81ff0658",
  1316 => x"5859758a",
  1317 => x"2e983876",
  1318 => x"81ff0651",
  1319 => x"e0a63f81",
  1320 => x"18587978",
  1321 => x"24e13879",
  1322 => x"b00c8d3d",
  1323 => x"0d048d51",
  1324 => x"e0923f78",
  1325 => x"337081ff",
  1326 => x"065257e0",
  1327 => x"873f8118",
  1328 => x"58e03979",
  1329 => x"557a547d",
  1330 => x"5385528d",
  1331 => x"3dfc0551",
  1332 => x"deef3fb0",
  1333 => x"0856868b",
  1334 => x"3f7bb008",
  1335 => x"0c75b00c",
  1336 => x"8d3d0d04",
  1337 => x"f63d0d7d",
  1338 => x"7f80c888",
  1339 => x"08705b58",
  1340 => x"5a5a7580",
  1341 => x"c1387779",
  1342 => x"25b338df",
  1343 => x"a23fb008",
  1344 => x"81ff0670",
  1345 => x"8d327030",
  1346 => x"709f2a51",
  1347 => x"51575776",
  1348 => x"8a2e80c3",
  1349 => x"3875802e",
  1350 => x"be38771a",
  1351 => x"56767634",
  1352 => x"7651dfa0",
  1353 => x"3f811858",
  1354 => x"787824cf",
  1355 => x"38775675",
  1356 => x"b00c8c3d",
  1357 => x"0d047855",
  1358 => x"79547c53",
  1359 => x"84528c3d",
  1360 => x"fc0551dd",
  1361 => x"fc3fb008",
  1362 => x"5685983f",
  1363 => x"7ab0080c",
  1364 => x"75b00c8c",
  1365 => x"3d0d0477",
  1366 => x"1a568a76",
  1367 => x"34811858",
  1368 => x"8d51dee0",
  1369 => x"3f8a51de",
  1370 => x"db3f7756",
  1371 => x"c239f93d",
  1372 => x"0d795780",
  1373 => x"c8880880",
  1374 => x"2eac3876",
  1375 => x"51879b3f",
  1376 => x"7b567a55",
  1377 => x"b0088105",
  1378 => x"54765382",
  1379 => x"52893dfc",
  1380 => x"0551ddad",
  1381 => x"3fb00857",
  1382 => x"84c93f77",
  1383 => x"b0080c76",
  1384 => x"b00c893d",
  1385 => x"0d0484bb",
  1386 => x"3f850bb0",
  1387 => x"080cff0b",
  1388 => x"b00c893d",
  1389 => x"0d04fb3d",
  1390 => x"0d80c888",
  1391 => x"08705654",
  1392 => x"73883874",
  1393 => x"b00c873d",
  1394 => x"0d047753",
  1395 => x"8352873d",
  1396 => x"fc0551dc",
  1397 => x"ec3fb008",
  1398 => x"5484883f",
  1399 => x"75b0080c",
  1400 => x"73b00c87",
  1401 => x"3d0d04ff",
  1402 => x"0bb00c04",
  1403 => x"fb3d0d77",
  1404 => x"5580c888",
  1405 => x"08802ea8",
  1406 => x"38745186",
  1407 => x"9d3fb008",
  1408 => x"81055474",
  1409 => x"53875287",
  1410 => x"3dfc0551",
  1411 => x"dcb33fb0",
  1412 => x"085583cf",
  1413 => x"3f75b008",
  1414 => x"0c74b00c",
  1415 => x"873d0d04",
  1416 => x"83c13f85",
  1417 => x"0bb0080c",
  1418 => x"ff0bb00c",
  1419 => x"873d0d04",
  1420 => x"fa3d0d80",
  1421 => x"c8880880",
  1422 => x"2ea2387a",
  1423 => x"55795478",
  1424 => x"53865288",
  1425 => x"3dfc0551",
  1426 => x"dbf73fb0",
  1427 => x"08568393",
  1428 => x"3f76b008",
  1429 => x"0c75b00c",
  1430 => x"883d0d04",
  1431 => x"83853f9d",
  1432 => x"0bb0080c",
  1433 => x"ff0bb00c",
  1434 => x"883d0d04",
  1435 => x"fb3d0d77",
  1436 => x"79565680",
  1437 => x"70545473",
  1438 => x"75259f38",
  1439 => x"74101010",
  1440 => x"f8055272",
  1441 => x"16703370",
  1442 => x"742b7607",
  1443 => x"8116f816",
  1444 => x"56565651",
  1445 => x"51747324",
  1446 => x"ea3873b0",
  1447 => x"0c873d0d",
  1448 => x"04fc3d0d",
  1449 => x"76785555",
  1450 => x"bc538052",
  1451 => x"735183db",
  1452 => x"3f845274",
  1453 => x"51ffb53f",
  1454 => x"b0087423",
  1455 => x"84528415",
  1456 => x"51ffa93f",
  1457 => x"b0088215",
  1458 => x"23845288",
  1459 => x"1551ff9c",
  1460 => x"3fb00884",
  1461 => x"150c8452",
  1462 => x"8c1551ff",
  1463 => x"8f3fb008",
  1464 => x"88152384",
  1465 => x"52901551",
  1466 => x"ff823fb0",
  1467 => x"088a1523",
  1468 => x"84529415",
  1469 => x"51fef53f",
  1470 => x"b0088c15",
  1471 => x"23845298",
  1472 => x"1551fee8",
  1473 => x"3fb0088e",
  1474 => x"15238852",
  1475 => x"9c1551fe",
  1476 => x"db3fb008",
  1477 => x"90150c86",
  1478 => x"3d0d04e9",
  1479 => x"3d0d6a80",
  1480 => x"c8880857",
  1481 => x"57759338",
  1482 => x"80c0800b",
  1483 => x"84180c75",
  1484 => x"ac180c75",
  1485 => x"b00c993d",
  1486 => x"0d04893d",
  1487 => x"70556a54",
  1488 => x"558a5299",
  1489 => x"3dffbc05",
  1490 => x"51d9f63f",
  1491 => x"b0087753",
  1492 => x"755256fe",
  1493 => x"cc3f818b",
  1494 => x"3f77b008",
  1495 => x"0c75b00c",
  1496 => x"993d0d04",
  1497 => x"e93d0d69",
  1498 => x"5780c888",
  1499 => x"08802eb5",
  1500 => x"38765183",
  1501 => x"a53f893d",
  1502 => x"7056b008",
  1503 => x"81055577",
  1504 => x"54568f52",
  1505 => x"993dffbc",
  1506 => x"0551d9b5",
  1507 => x"3fb0086b",
  1508 => x"53765257",
  1509 => x"fe8b3f80",
  1510 => x"ca3f77b0",
  1511 => x"080c76b0",
  1512 => x"0c993d0d",
  1513 => x"04bd3f85",
  1514 => x"0bb0080c",
  1515 => x"ff0bb00c",
  1516 => x"993d0d04",
  1517 => x"fc3d0d81",
  1518 => x"5480c888",
  1519 => x"08883873",
  1520 => x"b00c863d",
  1521 => x"0d047653",
  1522 => x"97b95286",
  1523 => x"3dfc0551",
  1524 => x"d8ef3fb0",
  1525 => x"08548c3f",
  1526 => x"74b0080c",
  1527 => x"73b00c86",
  1528 => x"3d0d04bf",
  1529 => x"d408b00c",
  1530 => x"04f73d0d",
  1531 => x"7bbfd408",
  1532 => x"82c81108",
  1533 => x"5a545a77",
  1534 => x"802e80d9",
  1535 => x"38818818",
  1536 => x"841908ff",
  1537 => x"0581712b",
  1538 => x"59555980",
  1539 => x"742480e9",
  1540 => x"38807424",
  1541 => x"b5387382",
  1542 => x"2b781188",
  1543 => x"05565681",
  1544 => x"80190877",
  1545 => x"06537280",
  1546 => x"2eb53878",
  1547 => x"16700853",
  1548 => x"53795174",
  1549 => x"0853722d",
  1550 => x"ff14fc17",
  1551 => x"fc177981",
  1552 => x"2c5a5757",
  1553 => x"54738025",
  1554 => x"d6387708",
  1555 => x"5877ffad",
  1556 => x"38bfd408",
  1557 => x"53bc1308",
  1558 => x"a5387951",
  1559 => x"f88c3f74",
  1560 => x"0853722d",
  1561 => x"ff14fc17",
  1562 => x"fc177981",
  1563 => x"2c5a5757",
  1564 => x"54738025",
  1565 => x"ffa938d2",
  1566 => x"398057ff",
  1567 => x"94397251",
  1568 => x"bc130853",
  1569 => x"722d7951",
  1570 => x"f7e03ffc",
  1571 => x"3d0d7679",
  1572 => x"71028c05",
  1573 => x"9f053357",
  1574 => x"55535583",
  1575 => x"72278a38",
  1576 => x"74830651",
  1577 => x"70802ea2",
  1578 => x"38ff1252",
  1579 => x"71ff2e93",
  1580 => x"38737370",
  1581 => x"81055534",
  1582 => x"ff125271",
  1583 => x"ff2e0981",
  1584 => x"06ef3874",
  1585 => x"b00c863d",
  1586 => x"0d047474",
  1587 => x"882b7507",
  1588 => x"7071902b",
  1589 => x"07515451",
  1590 => x"8f7227a5",
  1591 => x"38727170",
  1592 => x"8405530c",
  1593 => x"72717084",
  1594 => x"05530c72",
  1595 => x"71708405",
  1596 => x"530c7271",
  1597 => x"70840553",
  1598 => x"0cf01252",
  1599 => x"718f26dd",
  1600 => x"38837227",
  1601 => x"90387271",
  1602 => x"70840553",
  1603 => x"0cfc1252",
  1604 => x"718326f2",
  1605 => x"387053ff",
  1606 => x"9039fd3d",
  1607 => x"0d757071",
  1608 => x"83065355",
  1609 => x"5270b838",
  1610 => x"71700870",
  1611 => x"09f7fbfd",
  1612 => x"ff120670",
  1613 => x"f8848281",
  1614 => x"80065151",
  1615 => x"5253709d",
  1616 => x"38841370",
  1617 => x"087009f7",
  1618 => x"fbfdff12",
  1619 => x"0670f884",
  1620 => x"82818006",
  1621 => x"51515253",
  1622 => x"70802ee5",
  1623 => x"38725271",
  1624 => x"33517080",
  1625 => x"2e8a3881",
  1626 => x"12703352",
  1627 => x"5270f838",
  1628 => x"717431b0",
  1629 => x"0c853d0d",
  1630 => x"04ff3d0d",
  1631 => x"80c6d80b",
  1632 => x"fc057008",
  1633 => x"525270ff",
  1634 => x"2e913870",
  1635 => x"2dfc1270",
  1636 => x"08525270",
  1637 => x"ff2e0981",
  1638 => x"06f13883",
  1639 => x"3d0d0404",
  1640 => x"d8893f04",
  1641 => x"00ffffff",
  1642 => x"ff00ffff",
  1643 => x"ffff00ff",
  1644 => x"ffffff00",
  1645 => x"00000040",
  1646 => x"44485259",
  1647 => x"53544f4e",
  1648 => x"45205052",
  1649 => x"4f475241",
  1650 => x"4d2c2053",
  1651 => x"4f4d4520",
  1652 => x"53545249",
  1653 => x"4e470000",
  1654 => x"44485259",
  1655 => x"53544f4e",
  1656 => x"45205052",
  1657 => x"4f475241",
  1658 => x"4d2c2031",
  1659 => x"27535420",
  1660 => x"53545249",
  1661 => x"4e470000",
  1662 => x"44687279",
  1663 => x"73746f6e",
  1664 => x"65204265",
  1665 => x"6e63686d",
  1666 => x"61726b2c",
  1667 => x"20566572",
  1668 => x"73696f6e",
  1669 => x"20322e31",
  1670 => x"20284c61",
  1671 => x"6e677561",
  1672 => x"67653a20",
  1673 => x"43290a00",
  1674 => x"50726f67",
  1675 => x"72616d20",
  1676 => x"636f6d70",
  1677 => x"696c6564",
  1678 => x"20776974",
  1679 => x"68202772",
  1680 => x"65676973",
  1681 => x"74657227",
  1682 => x"20617474",
  1683 => x"72696275",
  1684 => x"74650a00",
  1685 => x"45786563",
  1686 => x"7574696f",
  1687 => x"6e207374",
  1688 => x"61727473",
  1689 => x"2c202564",
  1690 => x"2072756e",
  1691 => x"73207468",
  1692 => x"726f7567",
  1693 => x"68204468",
  1694 => x"72797374",
  1695 => x"6f6e650a",
  1696 => x"00000000",
  1697 => x"44485259",
  1698 => x"53544f4e",
  1699 => x"45205052",
  1700 => x"4f475241",
  1701 => x"4d2c2032",
  1702 => x"274e4420",
  1703 => x"53545249",
  1704 => x"4e470000",
  1705 => x"45786563",
  1706 => x"7574696f",
  1707 => x"6e20656e",
  1708 => x"64730a00",
  1709 => x"46696e61",
  1710 => x"6c207661",
  1711 => x"6c756573",
  1712 => x"206f6620",
  1713 => x"74686520",
  1714 => x"76617269",
  1715 => x"61626c65",
  1716 => x"73207573",
  1717 => x"65642069",
  1718 => x"6e207468",
  1719 => x"65206265",
  1720 => x"6e63686d",
  1721 => x"61726b3a",
  1722 => x"0a000000",
  1723 => x"496e745f",
  1724 => x"476c6f62",
  1725 => x"3a202020",
  1726 => x"20202020",
  1727 => x"20202020",
  1728 => x"2025640a",
  1729 => x"00000000",
  1730 => x"20202020",
  1731 => x"20202020",
  1732 => x"73686f75",
  1733 => x"6c642062",
  1734 => x"653a2020",
  1735 => x"2025640a",
  1736 => x"00000000",
  1737 => x"426f6f6c",
  1738 => x"5f476c6f",
  1739 => x"623a2020",
  1740 => x"20202020",
  1741 => x"20202020",
  1742 => x"2025640a",
  1743 => x"00000000",
  1744 => x"43685f31",
  1745 => x"5f476c6f",
  1746 => x"623a2020",
  1747 => x"20202020",
  1748 => x"20202020",
  1749 => x"2025630a",
  1750 => x"00000000",
  1751 => x"20202020",
  1752 => x"20202020",
  1753 => x"73686f75",
  1754 => x"6c642062",
  1755 => x"653a2020",
  1756 => x"2025630a",
  1757 => x"00000000",
  1758 => x"43685f32",
  1759 => x"5f476c6f",
  1760 => x"623a2020",
  1761 => x"20202020",
  1762 => x"20202020",
  1763 => x"2025630a",
  1764 => x"00000000",
  1765 => x"4172725f",
  1766 => x"315f476c",
  1767 => x"6f625b38",
  1768 => x"5d3a2020",
  1769 => x"20202020",
  1770 => x"2025640a",
  1771 => x"00000000",
  1772 => x"4172725f",
  1773 => x"325f476c",
  1774 => x"6f625b38",
  1775 => x"5d5b375d",
  1776 => x"3a202020",
  1777 => x"2025640a",
  1778 => x"00000000",
  1779 => x"20202020",
  1780 => x"20202020",
  1781 => x"73686f75",
  1782 => x"6c642062",
  1783 => x"653a2020",
  1784 => x"204e756d",
  1785 => x"6265725f",
  1786 => x"4f665f52",
  1787 => x"756e7320",
  1788 => x"2b203130",
  1789 => x"0a000000",
  1790 => x"5074725f",
  1791 => x"476c6f62",
  1792 => x"2d3e0a00",
  1793 => x"20205074",
  1794 => x"725f436f",
  1795 => x"6d703a20",
  1796 => x"20202020",
  1797 => x"20202020",
  1798 => x"2025640a",
  1799 => x"00000000",
  1800 => x"20202020",
  1801 => x"20202020",
  1802 => x"73686f75",
  1803 => x"6c642062",
  1804 => x"653a2020",
  1805 => x"2028696d",
  1806 => x"706c656d",
  1807 => x"656e7461",
  1808 => x"74696f6e",
  1809 => x"2d646570",
  1810 => x"656e6465",
  1811 => x"6e74290a",
  1812 => x"00000000",
  1813 => x"20204469",
  1814 => x"7363723a",
  1815 => x"20202020",
  1816 => x"20202020",
  1817 => x"20202020",
  1818 => x"2025640a",
  1819 => x"00000000",
  1820 => x"2020456e",
  1821 => x"756d5f43",
  1822 => x"6f6d703a",
  1823 => x"20202020",
  1824 => x"20202020",
  1825 => x"2025640a",
  1826 => x"00000000",
  1827 => x"2020496e",
  1828 => x"745f436f",
  1829 => x"6d703a20",
  1830 => x"20202020",
  1831 => x"20202020",
  1832 => x"2025640a",
  1833 => x"00000000",
  1834 => x"20205374",
  1835 => x"725f436f",
  1836 => x"6d703a20",
  1837 => x"20202020",
  1838 => x"20202020",
  1839 => x"2025730a",
  1840 => x"00000000",
  1841 => x"20202020",
  1842 => x"20202020",
  1843 => x"73686f75",
  1844 => x"6c642062",
  1845 => x"653a2020",
  1846 => x"20444852",
  1847 => x"5953544f",
  1848 => x"4e452050",
  1849 => x"524f4752",
  1850 => x"414d2c20",
  1851 => x"534f4d45",
  1852 => x"20535452",
  1853 => x"494e470a",
  1854 => x"00000000",
  1855 => x"4e657874",
  1856 => x"5f507472",
  1857 => x"5f476c6f",
  1858 => x"622d3e0a",
  1859 => x"00000000",
  1860 => x"20202020",
  1861 => x"20202020",
  1862 => x"73686f75",
  1863 => x"6c642062",
  1864 => x"653a2020",
  1865 => x"2028696d",
  1866 => x"706c656d",
  1867 => x"656e7461",
  1868 => x"74696f6e",
  1869 => x"2d646570",
  1870 => x"656e6465",
  1871 => x"6e74292c",
  1872 => x"2073616d",
  1873 => x"65206173",
  1874 => x"2061626f",
  1875 => x"76650a00",
  1876 => x"496e745f",
  1877 => x"315f4c6f",
  1878 => x"633a2020",
  1879 => x"20202020",
  1880 => x"20202020",
  1881 => x"2025640a",
  1882 => x"00000000",
  1883 => x"496e745f",
  1884 => x"325f4c6f",
  1885 => x"633a2020",
  1886 => x"20202020",
  1887 => x"20202020",
  1888 => x"2025640a",
  1889 => x"00000000",
  1890 => x"496e745f",
  1891 => x"335f4c6f",
  1892 => x"633a2020",
  1893 => x"20202020",
  1894 => x"20202020",
  1895 => x"2025640a",
  1896 => x"00000000",
  1897 => x"456e756d",
  1898 => x"5f4c6f63",
  1899 => x"3a202020",
  1900 => x"20202020",
  1901 => x"20202020",
  1902 => x"2025640a",
  1903 => x"00000000",
  1904 => x"5374725f",
  1905 => x"315f4c6f",
  1906 => x"633a2020",
  1907 => x"20202020",
  1908 => x"20202020",
  1909 => x"2025730a",
  1910 => x"00000000",
  1911 => x"20202020",
  1912 => x"20202020",
  1913 => x"73686f75",
  1914 => x"6c642062",
  1915 => x"653a2020",
  1916 => x"20444852",
  1917 => x"5953544f",
  1918 => x"4e452050",
  1919 => x"524f4752",
  1920 => x"414d2c20",
  1921 => x"31275354",
  1922 => x"20535452",
  1923 => x"494e470a",
  1924 => x"00000000",
  1925 => x"5374725f",
  1926 => x"325f4c6f",
  1927 => x"633a2020",
  1928 => x"20202020",
  1929 => x"20202020",
  1930 => x"2025730a",
  1931 => x"00000000",
  1932 => x"20202020",
  1933 => x"20202020",
  1934 => x"73686f75",
  1935 => x"6c642062",
  1936 => x"653a2020",
  1937 => x"20444852",
  1938 => x"5953544f",
  1939 => x"4e452050",
  1940 => x"524f4752",
  1941 => x"414d2c20",
  1942 => x"32274e44",
  1943 => x"20535452",
  1944 => x"494e470a",
  1945 => x"00000000",
  1946 => x"55736572",
  1947 => x"2074696d",
  1948 => x"653a2025",
  1949 => x"640a0000",
  1950 => x"4d696372",
  1951 => x"6f736563",
  1952 => x"6f6e6473",
  1953 => x"20666f72",
  1954 => x"206f6e65",
  1955 => x"2072756e",
  1956 => x"20746872",
  1957 => x"6f756768",
  1958 => x"20446872",
  1959 => x"7973746f",
  1960 => x"6e653a20",
  1961 => x"00000000",
  1962 => x"2564200a",
  1963 => x"00000000",
  1964 => x"44687279",
  1965 => x"73746f6e",
  1966 => x"65732070",
  1967 => x"65722053",
  1968 => x"65636f6e",
  1969 => x"643a2020",
  1970 => x"20202020",
  1971 => x"20202020",
  1972 => x"20202020",
  1973 => x"20202020",
  1974 => x"20202020",
  1975 => x"00000000",
  1976 => x"56415820",
  1977 => x"4d495053",
  1978 => x"20726174",
  1979 => x"696e6720",
  1980 => x"2a203130",
  1981 => x"3030203d",
  1982 => x"20256420",
  1983 => x"0a000000",
  1984 => x"50726f67",
  1985 => x"72616d20",
  1986 => x"636f6d70",
  1987 => x"696c6564",
  1988 => x"20776974",
  1989 => x"686f7574",
  1990 => x"20277265",
  1991 => x"67697374",
  1992 => x"65722720",
  1993 => x"61747472",
  1994 => x"69627574",
  1995 => x"650a0000",
  1996 => x"4d656173",
  1997 => x"75726564",
  1998 => x"2074696d",
  1999 => x"6520746f",
  2000 => x"6f20736d",
  2001 => x"616c6c20",
  2002 => x"746f206f",
  2003 => x"62746169",
  2004 => x"6e206d65",
  2005 => x"616e696e",
  2006 => x"6766756c",
  2007 => x"20726573",
  2008 => x"756c7473",
  2009 => x"0a000000",
  2010 => x"506c6561",
  2011 => x"73652069",
  2012 => x"6e637265",
  2013 => x"61736520",
  2014 => x"6e756d62",
  2015 => x"6572206f",
  2016 => x"66207275",
  2017 => x"6e730a00",
  2018 => x"44485259",
  2019 => x"53544f4e",
  2020 => x"45205052",
  2021 => x"4f475241",
  2022 => x"4d2c2033",
  2023 => x"27524420",
  2024 => x"53545249",
  2025 => x"4e470000",
  2026 => x"64756d6d",
  2027 => x"792e6578",
  2028 => x"65000000",
  2029 => x"43000000",
  2030 => x"00000000",
  2031 => x"00000000",
  2032 => x"00000000",
  2033 => x"00002360",
  2034 => x"000061a8",
  2035 => x"00000000",
  2036 => x"00001fa8",
  2037 => x"00001fd8",
  2038 => x"00000000",
  2039 => x"00002240",
  2040 => x"0000229c",
  2041 => x"000022f8",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"00000000",
  2049 => x"00000000",
  2050 => x"00000000",
  2051 => x"00001fb4",
  2052 => x"00000000",
  2053 => x"00000000",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000001",
  2081 => x"330eabcd",
  2082 => x"1234e66d",
  2083 => x"deec0005",
  2084 => x"000b0000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000000",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"00000000",
  2209 => x"00000000",
  2210 => x"00000000",
  2211 => x"00000000",
  2212 => x"00000000",
  2213 => x"00000000",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"00000000",
  2217 => x"00000000",
  2218 => x"00000000",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000000",
  2244 => x"00000000",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"ffffffff",
  2262 => x"00000000",
  2263 => x"ffffffff",
  2264 => x"00000000",
  2265 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;


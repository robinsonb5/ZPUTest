-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_ROM;

architecture arch of Dhrystone_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"80700b0b",
     2 => x"80c0b00c",
     3 => x"3a0b0b0b",
     4 => x"a9810400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"8f040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bb4",
   162 => x"84738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f7040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"df040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80c0ac0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"83e13fab",
   257 => x"d23f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104b0",
   280 => x"08b408b8",
   281 => x"087575a3",
   282 => x"a72d5050",
   283 => x"b00856b8",
   284 => x"0cb40cb0",
   285 => x"0c5104b0",
   286 => x"08b408b8",
   287 => x"087575a1",
   288 => x"f52d5050",
   289 => x"b00856b8",
   290 => x"0cb40cb0",
   291 => x"0c5104b0",
   292 => x"08b408b8",
   293 => x"08a9c82d",
   294 => x"b80cb40c",
   295 => x"b00c04fe",
   296 => x"3d0d0b0b",
   297 => x"80c7dc08",
   298 => x"53841308",
   299 => x"70882a70",
   300 => x"81065152",
   301 => x"5270802e",
   302 => x"f0387181",
   303 => x"ff06b00c",
   304 => x"843d0d04",
   305 => x"ff3d0d0b",
   306 => x"0b80c7dc",
   307 => x"08527108",
   308 => x"70882a81",
   309 => x"32708106",
   310 => x"51515170",
   311 => x"f1387372",
   312 => x"0c833d0d",
   313 => x"0480c0ac",
   314 => x"08802ea4",
   315 => x"3880c0b0",
   316 => x"08822ebd",
   317 => x"38838080",
   318 => x"0b0b0b80",
   319 => x"c7dc0c82",
   320 => x"a0800b80",
   321 => x"c7e00c82",
   322 => x"90800b80",
   323 => x"c7e40c04",
   324 => x"f8808080",
   325 => x"a40b0b0b",
   326 => x"80c7dc0c",
   327 => x"f8808082",
   328 => x"800b80c7",
   329 => x"e00cf880",
   330 => x"8084800b",
   331 => x"80c7e40c",
   332 => x"0480c0a8",
   333 => x"808c0b0b",
   334 => x"0b80c7dc",
   335 => x"0c80c0a8",
   336 => x"80940b80",
   337 => x"c7e00cb4",
   338 => x"940b80c7",
   339 => x"e40c04f2",
   340 => x"3d0d6080",
   341 => x"c7e00856",
   342 => x"5d82750c",
   343 => x"8059805a",
   344 => x"800b8f3d",
   345 => x"5d5b7a10",
   346 => x"10157008",
   347 => x"7108719f",
   348 => x"2c7e852b",
   349 => x"5855557d",
   350 => x"53595795",
   351 => x"823f7d7f",
   352 => x"7a72077c",
   353 => x"72077171",
   354 => x"60810541",
   355 => x"5f5d5b59",
   356 => x"5755817b",
   357 => x"278f3876",
   358 => x"7d0c7784",
   359 => x"1e0c7cb0",
   360 => x"0c903d0d",
   361 => x"0480c7e0",
   362 => x"0855ffba",
   363 => x"39ff3d0d",
   364 => x"80c7e833",
   365 => x"5170a738",
   366 => x"80c0b808",
   367 => x"70085252",
   368 => x"70802e94",
   369 => x"38841280",
   370 => x"c0b80c70",
   371 => x"2d80c0b8",
   372 => x"08700852",
   373 => x"5270ee38",
   374 => x"810b80c7",
   375 => x"e834833d",
   376 => x"0d040480",
   377 => x"3d0d0b0b",
   378 => x"80c7d808",
   379 => x"802e8e38",
   380 => x"0b0b0b0b",
   381 => x"800b802e",
   382 => x"09810685",
   383 => x"38823d0d",
   384 => x"040b0b80",
   385 => x"c7d8510b",
   386 => x"0b0bf3f4",
   387 => x"3f823d0d",
   388 => x"0404c008",
   389 => x"b00c0480",
   390 => x"3d0d80c1",
   391 => x"0b8197cc",
   392 => x"34800b81",
   393 => x"99e40c70",
   394 => x"b00c823d",
   395 => x"0d04ff3d",
   396 => x"0d800b81",
   397 => x"97cc3352",
   398 => x"527080c1",
   399 => x"2e993871",
   400 => x"8199e408",
   401 => x"078199e4",
   402 => x"0c80c20b",
   403 => x"8197d034",
   404 => x"70b00c83",
   405 => x"3d0d0481",
   406 => x"0b8199e4",
   407 => x"08078199",
   408 => x"e40c80c2",
   409 => x"0b8197d0",
   410 => x"3470b00c",
   411 => x"833d0d04",
   412 => x"fd3d0d75",
   413 => x"70088a05",
   414 => x"53538197",
   415 => x"cc335170",
   416 => x"80c12e8b",
   417 => x"3873f338",
   418 => x"70b00c85",
   419 => x"3d0d04ff",
   420 => x"12708197",
   421 => x"c8083174",
   422 => x"0cb00c85",
   423 => x"3d0d04fc",
   424 => x"3d0d8197",
   425 => x"f4085574",
   426 => x"802e8c38",
   427 => x"76750871",
   428 => x"0c8197f4",
   429 => x"0856548c",
   430 => x"15538197",
   431 => x"c808528a",
   432 => x"518ca33f",
   433 => x"73b00c86",
   434 => x"3d0d04fb",
   435 => x"3d0d7770",
   436 => x"085656b0",
   437 => x"538197f4",
   438 => x"08527451",
   439 => x"98f53f85",
   440 => x"0b8c170c",
   441 => x"850b8c16",
   442 => x"0c750875",
   443 => x"0c8197f4",
   444 => x"08547380",
   445 => x"2e8a3873",
   446 => x"08750c81",
   447 => x"97f40854",
   448 => x"8c145381",
   449 => x"97c80852",
   450 => x"8a518bda",
   451 => x"3f841508",
   452 => x"ad38860b",
   453 => x"8c160c88",
   454 => x"15528816",
   455 => x"08518ae6",
   456 => x"3f8197f4",
   457 => x"08700876",
   458 => x"0c548c15",
   459 => x"7054548a",
   460 => x"52730851",
   461 => x"8bb03f73",
   462 => x"b00c873d",
   463 => x"0d047508",
   464 => x"54b05373",
   465 => x"52755198",
   466 => x"8a3f73b0",
   467 => x"0c873d0d",
   468 => x"04f33d0d",
   469 => x"88bd0bff",
   470 => x"880c8196",
   471 => x"e00b8197",
   472 => x"940c8197",
   473 => x"980b8197",
   474 => x"f40c8196",
   475 => x"e00b8197",
   476 => x"980c800b",
   477 => x"8197980b",
   478 => x"84050c82",
   479 => x"0b819798",
   480 => x"0b88050c",
   481 => x"a80b8197",
   482 => x"980b8c05",
   483 => x"0c9f53b4",
   484 => x"98528197",
   485 => x"a85197bb",
   486 => x"3f9f53b4",
   487 => x"b8528199",
   488 => x"c45197af",
   489 => x"3f8a0b80",
   490 => x"d5ac0cbe",
   491 => x"dc518dda",
   492 => x"3fb4d851",
   493 => x"8dd43fbe",
   494 => x"dc518dce",
   495 => x"3f80c0c0",
   496 => x"08802e87",
   497 => x"d238b588",
   498 => x"518dbf3f",
   499 => x"bedc518d",
   500 => x"b93f80c0",
   501 => x"bc0852b5",
   502 => x"b4518dae",
   503 => x"3fc00880",
   504 => x"c8cc0c81",
   505 => x"58800b80",
   506 => x"c0bc0825",
   507 => x"82d0388c",
   508 => x"3d5b80c1",
   509 => x"0b8197cc",
   510 => x"34810b81",
   511 => x"99e40c80",
   512 => x"c20b8197",
   513 => x"d034825c",
   514 => x"835a9f53",
   515 => x"b5e45281",
   516 => x"97d45196",
   517 => x"be3f815d",
   518 => x"800b8197",
   519 => x"d4538199",
   520 => x"c452558a",
   521 => x"e53fb008",
   522 => x"752e0981",
   523 => x"06833881",
   524 => x"55748199",
   525 => x"e40c7b70",
   526 => x"57557483",
   527 => x"25a03874",
   528 => x"101015fd",
   529 => x"055e8f3d",
   530 => x"fc055383",
   531 => x"52755189",
   532 => x"953f811c",
   533 => x"705d7057",
   534 => x"55837524",
   535 => x"e2387d54",
   536 => x"745380c8",
   537 => x"d0528197",
   538 => x"fc51898a",
   539 => x"3f8197f4",
   540 => x"08700857",
   541 => x"57b05376",
   542 => x"52755195",
   543 => x"d63f850b",
   544 => x"8c180c85",
   545 => x"0b8c170c",
   546 => x"7608760c",
   547 => x"8197f408",
   548 => x"5574802e",
   549 => x"8a387408",
   550 => x"760c8197",
   551 => x"f408558c",
   552 => x"15538197",
   553 => x"c808528a",
   554 => x"5188bb3f",
   555 => x"84160887",
   556 => x"8e38860b",
   557 => x"8c170c88",
   558 => x"16528817",
   559 => x"085187c6",
   560 => x"3f8197f4",
   561 => x"08700877",
   562 => x"0c558c16",
   563 => x"7054578a",
   564 => x"52760851",
   565 => x"88903f80",
   566 => x"c10b8197",
   567 => x"d0335656",
   568 => x"757526a2",
   569 => x"3880c352",
   570 => x"755188f4",
   571 => x"3fb0087d",
   572 => x"2e869f38",
   573 => x"81167081",
   574 => x"ff068197",
   575 => x"d0335757",
   576 => x"57747627",
   577 => x"e038797c",
   578 => x"297e7072",
   579 => x"35705f72",
   580 => x"72317087",
   581 => x"29723153",
   582 => x"538a0581",
   583 => x"97cc3381",
   584 => x"97c8085a",
   585 => x"5a525b55",
   586 => x"7680c12e",
   587 => x"86a93878",
   588 => x"f7388118",
   589 => x"5880c0bc",
   590 => x"087825fd",
   591 => x"b538c008",
   592 => x"8197900c",
   593 => x"b684518a",
   594 => x"c13fbedc",
   595 => x"518abb3f",
   596 => x"b694518a",
   597 => x"b53fbedc",
   598 => x"518aaf3f",
   599 => x"8197c808",
   600 => x"52b6cc51",
   601 => x"8aa43f85",
   602 => x"52b6e851",
   603 => x"8a9c3f81",
   604 => x"99e40852",
   605 => x"b784518a",
   606 => x"913f8152",
   607 => x"b6e8518a",
   608 => x"893f8197",
   609 => x"cc3352b7",
   610 => x"a05189fe",
   611 => x"3f80c152",
   612 => x"b7bc5189",
   613 => x"f53f8197",
   614 => x"d03352b7",
   615 => x"d85189ea",
   616 => x"3f80c252",
   617 => x"b7bc5189",
   618 => x"e13f8198",
   619 => x"9c0852b7",
   620 => x"f45189d6",
   621 => x"3f8752b6",
   622 => x"e85189ce",
   623 => x"3f80d5ac",
   624 => x"0852b890",
   625 => x"5189c33f",
   626 => x"b8ac5189",
   627 => x"bd3fb8d8",
   628 => x"5189b73f",
   629 => x"8197f408",
   630 => x"70085357",
   631 => x"b8e45189",
   632 => x"a93fb980",
   633 => x"5189a33f",
   634 => x"8197f408",
   635 => x"84110853",
   636 => x"5bb9b451",
   637 => x"89943f80",
   638 => x"52b6e851",
   639 => x"898c3f81",
   640 => x"97f40888",
   641 => x"11085358",
   642 => x"b9d05188",
   643 => x"fd3f8252",
   644 => x"b6e85188",
   645 => x"f53f8197",
   646 => x"f4088c11",
   647 => x"085359b9",
   648 => x"ec5188e6",
   649 => x"3f9152b6",
   650 => x"e85188de",
   651 => x"3f8197f4",
   652 => x"08900552",
   653 => x"ba885188",
   654 => x"d13fbaa4",
   655 => x"5188cb3f",
   656 => x"badc5188",
   657 => x"c53f8197",
   658 => x"94087008",
   659 => x"5355b8e4",
   660 => x"5188b73f",
   661 => x"baf05188",
   662 => x"b13f8197",
   663 => x"94088411",
   664 => x"085356b9",
   665 => x"b45188a2",
   666 => x"3f8052b6",
   667 => x"e851889a",
   668 => x"3f819794",
   669 => x"08881108",
   670 => x"5357b9d0",
   671 => x"51888b3f",
   672 => x"8152b6e8",
   673 => x"5188833f",
   674 => x"81979408",
   675 => x"8c110853",
   676 => x"5bb9ec51",
   677 => x"87f43f92",
   678 => x"52b6e851",
   679 => x"87ec3f81",
   680 => x"97940890",
   681 => x"0552ba88",
   682 => x"5187df3f",
   683 => x"baa45187",
   684 => x"d93f7b52",
   685 => x"bbb05187",
   686 => x"d13f8552",
   687 => x"b6e85187",
   688 => x"c93f7952",
   689 => x"bbcc5187",
   690 => x"c13f8d52",
   691 => x"b6e85187",
   692 => x"b93f7d52",
   693 => x"bbe85187",
   694 => x"b13f8752",
   695 => x"b6e85187",
   696 => x"a93f7c52",
   697 => x"bc845187",
   698 => x"a13f8152",
   699 => x"b6e85187",
   700 => x"993f8199",
   701 => x"c452bca0",
   702 => x"51878f3f",
   703 => x"bcbc5187",
   704 => x"893f8197",
   705 => x"d452bcf4",
   706 => x"5186ff3f",
   707 => x"bd905186",
   708 => x"f93fbedc",
   709 => x"5186f33f",
   710 => x"81979008",
   711 => x"80c8cc08",
   712 => x"317080c8",
   713 => x"c80c52bd",
   714 => x"c85186de",
   715 => x"3f80c8c8",
   716 => x"085680f7",
   717 => x"762580e5",
   718 => x"3880c0bc",
   719 => x"08707787",
   720 => x"e8293580",
   721 => x"c8c00c76",
   722 => x"7187e829",
   723 => x"3580c8c4",
   724 => x"0c767184",
   725 => x"b9293581",
   726 => x"97f80c5a",
   727 => x"bdd85186",
   728 => x"a93f80c8",
   729 => x"c00852be",
   730 => x"8851869e",
   731 => x"3fbe9051",
   732 => x"86983f80",
   733 => x"c8c40852",
   734 => x"be885186",
   735 => x"8d3f8197",
   736 => x"f80852be",
   737 => x"c0518682",
   738 => x"3fbedc51",
   739 => x"85fc3f80",
   740 => x"0bb00c8f",
   741 => x"3d0d04be",
   742 => x"e051f8ad",
   743 => x"39bf9051",
   744 => x"85e83fbf",
   745 => x"c85185e2",
   746 => x"3fbedc51",
   747 => x"85dc3f80",
   748 => x"c8c80880",
   749 => x"c0bc0870",
   750 => x"7287e829",
   751 => x"3580c8c0",
   752 => x"0c717187",
   753 => x"e8293580",
   754 => x"c8c40c71",
   755 => x"7184b929",
   756 => x"358197f8",
   757 => x"0c5b56bd",
   758 => x"d85185ae",
   759 => x"3f80c8c0",
   760 => x"0852be88",
   761 => x"5185a33f",
   762 => x"be905185",
   763 => x"9d3f80c8",
   764 => x"c40852be",
   765 => x"88518592",
   766 => x"3f8197f8",
   767 => x"0852bec0",
   768 => x"5185873f",
   769 => x"bedc5185",
   770 => x"813f800b",
   771 => x"b00c8f3d",
   772 => x"0d048f3d",
   773 => x"f8055280",
   774 => x"5180eb3f",
   775 => x"9f53bfe8",
   776 => x"528197d4",
   777 => x"518eac3f",
   778 => x"77788197",
   779 => x"c80c8117",
   780 => x"7081ff06",
   781 => x"8197d033",
   782 => x"5858585a",
   783 => x"f9c33976",
   784 => x"0856b053",
   785 => x"75527651",
   786 => x"8e893f80",
   787 => x"c10b8197",
   788 => x"d0335656",
   789 => x"f98a39ff",
   790 => x"15707731",
   791 => x"7c0c5980",
   792 => x"0b811959",
   793 => x"5980c0bc",
   794 => x"087825f7",
   795 => x"8538f9ce",
   796 => x"39ff3d0d",
   797 => x"73823270",
   798 => x"30707207",
   799 => x"8025b00c",
   800 => x"5252833d",
   801 => x"0d04fe3d",
   802 => x"0d747671",
   803 => x"53545271",
   804 => x"822e8338",
   805 => x"83517181",
   806 => x"2e9a3881",
   807 => x"72269f38",
   808 => x"71822eb8",
   809 => x"3871842e",
   810 => x"a9387073",
   811 => x"0c70b00c",
   812 => x"843d0d04",
   813 => x"80e40b81",
   814 => x"97c80825",
   815 => x"8b388073",
   816 => x"0c70b00c",
   817 => x"843d0d04",
   818 => x"83730c70",
   819 => x"b00c843d",
   820 => x"0d048273",
   821 => x"0c70b00c",
   822 => x"843d0d04",
   823 => x"81730c70",
   824 => x"b00c843d",
   825 => x"0d04803d",
   826 => x"0d747414",
   827 => x"8205710c",
   828 => x"b00c823d",
   829 => x"0d04f73d",
   830 => x"0d7b7d7f",
   831 => x"61851270",
   832 => x"822b7511",
   833 => x"70747170",
   834 => x"8405530c",
   835 => x"5a5a5d5b",
   836 => x"760c7980",
   837 => x"f8180c79",
   838 => x"86125257",
   839 => x"585a5a76",
   840 => x"76249938",
   841 => x"76b32982",
   842 => x"2b791151",
   843 => x"53767370",
   844 => x"8405550c",
   845 => x"81145475",
   846 => x"7425f238",
   847 => x"7681cc29",
   848 => x"19fc1108",
   849 => x"8105fc12",
   850 => x"0c7a1970",
   851 => x"089fa013",
   852 => x"0c585685",
   853 => x"0b8197c8",
   854 => x"0c75b00c",
   855 => x"8b3d0d04",
   856 => x"fe3d0d02",
   857 => x"93053351",
   858 => x"80028405",
   859 => x"97053354",
   860 => x"5270732e",
   861 => x"883871b0",
   862 => x"0c843d0d",
   863 => x"04708197",
   864 => x"cc34810b",
   865 => x"b00c843d",
   866 => x"0d04f83d",
   867 => x"0d7a7c59",
   868 => x"56820b83",
   869 => x"19555574",
   870 => x"16703375",
   871 => x"335b5153",
   872 => x"72792e80",
   873 => x"c63880c1",
   874 => x"0b811681",
   875 => x"16565657",
   876 => x"827525e3",
   877 => x"38ffa917",
   878 => x"7081ff06",
   879 => x"55597382",
   880 => x"26833887",
   881 => x"55815376",
   882 => x"80d22e98",
   883 => x"38775275",
   884 => x"518c993f",
   885 => x"805372b0",
   886 => x"08258938",
   887 => x"87158197",
   888 => x"c80c8153",
   889 => x"72b00c8a",
   890 => x"3d0d0472",
   891 => x"8197cc34",
   892 => x"827525ff",
   893 => x"a238ffbd",
   894 => x"39ff3d0d",
   895 => x"028f0533",
   896 => x"52ff8408",
   897 => x"70882a70",
   898 => x"81065151",
   899 => x"5170802e",
   900 => x"f03871ff",
   901 => x"840c833d",
   902 => x"0d04fe3d",
   903 => x"0d747033",
   904 => x"52537080",
   905 => x"2ea13870",
   906 => x"52811353",
   907 => x"ff840870",
   908 => x"882a7081",
   909 => x"06515151",
   910 => x"70802ef0",
   911 => x"3871ff84",
   912 => x"0c723352",
   913 => x"71e33884",
   914 => x"3d0d04ff",
   915 => x"3d0dff84",
   916 => x"0870892a",
   917 => x"70810651",
   918 => x"52527080",
   919 => x"2ef03871",
   920 => x"81ff06b0",
   921 => x"0c833d0d",
   922 => x"04ff3d0d",
   923 => x"028f0533",
   924 => x"52ff8408",
   925 => x"70882a70",
   926 => x"81065151",
   927 => x"5170802e",
   928 => x"f03871ff",
   929 => x"840c833d",
   930 => x"0d04f53d",
   931 => x"0d8e3d70",
   932 => x"70840552",
   933 => x"089ce95b",
   934 => x"555b8074",
   935 => x"70810556",
   936 => x"33755a54",
   937 => x"5772772e",
   938 => x"be3872a5",
   939 => x"2e098106",
   940 => x"80c53877",
   941 => x"70810559",
   942 => x"33537280",
   943 => x"e42e81b6",
   944 => x"387280e4",
   945 => x"2480c638",
   946 => x"7280e32e",
   947 => x"a1388052",
   948 => x"a551782d",
   949 => x"80527251",
   950 => x"782d8217",
   951 => x"57777081",
   952 => x"05593353",
   953 => x"72c43876",
   954 => x"b00c8d3d",
   955 => x"0d047a84",
   956 => x"1c831233",
   957 => x"555c5680",
   958 => x"52725178",
   959 => x"2d811778",
   960 => x"7081055a",
   961 => x"33545772",
   962 => x"ffa038db",
   963 => x"397280f3",
   964 => x"2e098106",
   965 => x"ffb8387a",
   966 => x"841c7108",
   967 => x"585c5480",
   968 => x"76335b55",
   969 => x"79752e8d",
   970 => x"38811570",
   971 => x"17703355",
   972 => x"5b5572f5",
   973 => x"38ff1554",
   974 => x"807525ff",
   975 => x"a0387570",
   976 => x"81055733",
   977 => x"53805272",
   978 => x"51782d81",
   979 => x"1774ff16",
   980 => x"56565780",
   981 => x"7525ff85",
   982 => x"38757081",
   983 => x"05573353",
   984 => x"80527251",
   985 => x"782d8117",
   986 => x"74ff1656",
   987 => x"56577480",
   988 => x"24cc38fe",
   989 => x"e8397a84",
   990 => x"1c710881",
   991 => x"99f80b80",
   992 => x"c7ec545d",
   993 => x"565c5580",
   994 => x"5673762e",
   995 => x"098106b8",
   996 => x"38b00b80",
   997 => x"c7ec3481",
   998 => x"1555ff15",
   999 => x"5574337a",
  1000 => x"7081055c",
  1001 => x"34811656",
  1002 => x"7480c7ec",
  1003 => x"2e098106",
  1004 => x"e938807a",
  1005 => x"34758199",
  1006 => x"f80bff12",
  1007 => x"56575574",
  1008 => x"8024fefa",
  1009 => x"38fe9639",
  1010 => x"738f0680",
  1011 => x"c0880553",
  1012 => x"72337570",
  1013 => x"81055734",
  1014 => x"73842a54",
  1015 => x"73ea3874",
  1016 => x"80c7ec2e",
  1017 => x"cd38ff15",
  1018 => x"5574337a",
  1019 => x"7081055c",
  1020 => x"34811656",
  1021 => x"7480c7ec",
  1022 => x"2effb738",
  1023 => x"ff9c39bc",
  1024 => x"0802bc0c",
  1025 => x"f53d0dbc",
  1026 => x"08940508",
  1027 => x"9d38bc08",
  1028 => x"8c0508bc",
  1029 => x"08900508",
  1030 => x"bc088805",
  1031 => x"08585654",
  1032 => x"73760c74",
  1033 => x"84170c81",
  1034 => x"bf39800b",
  1035 => x"bc08f005",
  1036 => x"0c800bbc",
  1037 => x"08f4050c",
  1038 => x"bc088c05",
  1039 => x"08bc0890",
  1040 => x"05085654",
  1041 => x"73bc08f0",
  1042 => x"050c74bc",
  1043 => x"08f4050c",
  1044 => x"bc08f805",
  1045 => x"bc08f005",
  1046 => x"56568870",
  1047 => x"54755376",
  1048 => x"525485ef",
  1049 => x"3fa00bbc",
  1050 => x"08940508",
  1051 => x"31bc08ec",
  1052 => x"050cbc08",
  1053 => x"ec050880",
  1054 => x"249d3880",
  1055 => x"0bbc08f4",
  1056 => x"050cbc08",
  1057 => x"ec050830",
  1058 => x"bc08fc05",
  1059 => x"08712bbc",
  1060 => x"08f0050c",
  1061 => x"54b939bc",
  1062 => x"08fc0508",
  1063 => x"bc08ec05",
  1064 => x"082abc08",
  1065 => x"e8050cbc",
  1066 => x"08fc0508",
  1067 => x"bc089405",
  1068 => x"082bbc08",
  1069 => x"f4050cbc",
  1070 => x"08f80508",
  1071 => x"bc089405",
  1072 => x"082b70bc",
  1073 => x"08e80508",
  1074 => x"07bc08f0",
  1075 => x"050c54bc",
  1076 => x"08f00508",
  1077 => x"bc08f405",
  1078 => x"08bc0888",
  1079 => x"05085856",
  1080 => x"5473760c",
  1081 => x"7484170c",
  1082 => x"bc088805",
  1083 => x"08b00c8d",
  1084 => x"3d0dbc0c",
  1085 => x"04bc0802",
  1086 => x"bc0cf93d",
  1087 => x"0d800bbc",
  1088 => x"08fc050c",
  1089 => x"bc088805",
  1090 => x"088025ab",
  1091 => x"38bc0888",
  1092 => x"050830bc",
  1093 => x"0888050c",
  1094 => x"800bbc08",
  1095 => x"f4050cbc",
  1096 => x"08fc0508",
  1097 => x"8838810b",
  1098 => x"bc08f405",
  1099 => x"0cbc08f4",
  1100 => x"0508bc08",
  1101 => x"fc050cbc",
  1102 => x"088c0508",
  1103 => x"8025ab38",
  1104 => x"bc088c05",
  1105 => x"0830bc08",
  1106 => x"8c050c80",
  1107 => x"0bbc08f0",
  1108 => x"050cbc08",
  1109 => x"fc050888",
  1110 => x"38810bbc",
  1111 => x"08f0050c",
  1112 => x"bc08f005",
  1113 => x"08bc08fc",
  1114 => x"050c8053",
  1115 => x"bc088c05",
  1116 => x"0852bc08",
  1117 => x"88050851",
  1118 => x"81a73fb0",
  1119 => x"0870bc08",
  1120 => x"f8050c54",
  1121 => x"bc08fc05",
  1122 => x"08802e8c",
  1123 => x"38bc08f8",
  1124 => x"050830bc",
  1125 => x"08f8050c",
  1126 => x"bc08f805",
  1127 => x"0870b00c",
  1128 => x"54893d0d",
  1129 => x"bc0c04bc",
  1130 => x"0802bc0c",
  1131 => x"fb3d0d80",
  1132 => x"0bbc08fc",
  1133 => x"050cbc08",
  1134 => x"88050880",
  1135 => x"259338bc",
  1136 => x"08880508",
  1137 => x"30bc0888",
  1138 => x"050c810b",
  1139 => x"bc08fc05",
  1140 => x"0cbc088c",
  1141 => x"05088025",
  1142 => x"8c38bc08",
  1143 => x"8c050830",
  1144 => x"bc088c05",
  1145 => x"0c8153bc",
  1146 => x"088c0508",
  1147 => x"52bc0888",
  1148 => x"050851ad",
  1149 => x"3fb00870",
  1150 => x"bc08f805",
  1151 => x"0c54bc08",
  1152 => x"fc050880",
  1153 => x"2e8c38bc",
  1154 => x"08f80508",
  1155 => x"30bc08f8",
  1156 => x"050cbc08",
  1157 => x"f8050870",
  1158 => x"b00c5487",
  1159 => x"3d0dbc0c",
  1160 => x"04bc0802",
  1161 => x"bc0cfd3d",
  1162 => x"0d810bbc",
  1163 => x"08fc050c",
  1164 => x"800bbc08",
  1165 => x"f8050cbc",
  1166 => x"088c0508",
  1167 => x"bc088805",
  1168 => x"0827ac38",
  1169 => x"bc08fc05",
  1170 => x"08802ea3",
  1171 => x"38800bbc",
  1172 => x"088c0508",
  1173 => x"249938bc",
  1174 => x"088c0508",
  1175 => x"10bc088c",
  1176 => x"050cbc08",
  1177 => x"fc050810",
  1178 => x"bc08fc05",
  1179 => x"0cc939bc",
  1180 => x"08fc0508",
  1181 => x"802e80c9",
  1182 => x"38bc088c",
  1183 => x"0508bc08",
  1184 => x"88050826",
  1185 => x"a138bc08",
  1186 => x"880508bc",
  1187 => x"088c0508",
  1188 => x"31bc0888",
  1189 => x"050cbc08",
  1190 => x"f80508bc",
  1191 => x"08fc0508",
  1192 => x"07bc08f8",
  1193 => x"050cbc08",
  1194 => x"fc050881",
  1195 => x"2abc08fc",
  1196 => x"050cbc08",
  1197 => x"8c050881",
  1198 => x"2abc088c",
  1199 => x"050cffaf",
  1200 => x"39bc0890",
  1201 => x"0508802e",
  1202 => x"8f38bc08",
  1203 => x"88050870",
  1204 => x"bc08f405",
  1205 => x"0c518d39",
  1206 => x"bc08f805",
  1207 => x"0870bc08",
  1208 => x"f4050c51",
  1209 => x"bc08f405",
  1210 => x"08b00c85",
  1211 => x"3d0dbc0c",
  1212 => x"04bc0802",
  1213 => x"bc0cff3d",
  1214 => x"0d800bbc",
  1215 => x"08fc050c",
  1216 => x"bc088805",
  1217 => x"088106ff",
  1218 => x"11700970",
  1219 => x"bc088c05",
  1220 => x"0806bc08",
  1221 => x"fc050811",
  1222 => x"bc08fc05",
  1223 => x"0cbc0888",
  1224 => x"0508812a",
  1225 => x"bc088805",
  1226 => x"0cbc088c",
  1227 => x"050810bc",
  1228 => x"088c050c",
  1229 => x"51515151",
  1230 => x"bc088805",
  1231 => x"08802e84",
  1232 => x"38ffbd39",
  1233 => x"bc08fc05",
  1234 => x"0870b00c",
  1235 => x"51833d0d",
  1236 => x"bc0c04fc",
  1237 => x"3d0d7670",
  1238 => x"797b5555",
  1239 => x"55558f72",
  1240 => x"278c3872",
  1241 => x"75078306",
  1242 => x"5170802e",
  1243 => x"a738ff12",
  1244 => x"5271ff2e",
  1245 => x"98387270",
  1246 => x"81055433",
  1247 => x"74708105",
  1248 => x"5634ff12",
  1249 => x"5271ff2e",
  1250 => x"098106ea",
  1251 => x"3874b00c",
  1252 => x"863d0d04",
  1253 => x"74517270",
  1254 => x"84055408",
  1255 => x"71708405",
  1256 => x"530c7270",
  1257 => x"84055408",
  1258 => x"71708405",
  1259 => x"530c7270",
  1260 => x"84055408",
  1261 => x"71708405",
  1262 => x"530c7270",
  1263 => x"84055408",
  1264 => x"71708405",
  1265 => x"530cf012",
  1266 => x"52718f26",
  1267 => x"c9388372",
  1268 => x"27953872",
  1269 => x"70840554",
  1270 => x"08717084",
  1271 => x"05530cfc",
  1272 => x"12527183",
  1273 => x"26ed3870",
  1274 => x"54ff8339",
  1275 => x"fb3d0d77",
  1276 => x"79707207",
  1277 => x"83065354",
  1278 => x"52709338",
  1279 => x"71737308",
  1280 => x"54565471",
  1281 => x"73082e80",
  1282 => x"c4387375",
  1283 => x"54527133",
  1284 => x"7081ff06",
  1285 => x"52547080",
  1286 => x"2e9d3872",
  1287 => x"33557075",
  1288 => x"2e098106",
  1289 => x"95388112",
  1290 => x"81147133",
  1291 => x"7081ff06",
  1292 => x"54565452",
  1293 => x"70e53872",
  1294 => x"33557381",
  1295 => x"ff067581",
  1296 => x"ff067171",
  1297 => x"31b00c52",
  1298 => x"52873d0d",
  1299 => x"04710970",
  1300 => x"f7fbfdff",
  1301 => x"140670f8",
  1302 => x"84828180",
  1303 => x"06515151",
  1304 => x"70973884",
  1305 => x"14841671",
  1306 => x"08545654",
  1307 => x"7175082e",
  1308 => x"dc387375",
  1309 => x"5452ff96",
  1310 => x"39800bb0",
  1311 => x"0c873d0d",
  1312 => x"04fd3d0d",
  1313 => x"800b80c0",
  1314 => x"b0085454",
  1315 => x"72812e9b",
  1316 => x"387380c8",
  1317 => x"bc0ce0cd",
  1318 => x"3fdee53f",
  1319 => x"80c0c452",
  1320 => x"8151e5ad",
  1321 => x"3fb00851",
  1322 => x"879b3f72",
  1323 => x"80c8bc0c",
  1324 => x"e0b33fde",
  1325 => x"cb3f80c0",
  1326 => x"c4528151",
  1327 => x"e5933fb0",
  1328 => x"08518781",
  1329 => x"3f00ff39",
  1330 => x"00ff39f5",
  1331 => x"3d0d7e60",
  1332 => x"80c8bc08",
  1333 => x"705b585b",
  1334 => x"5b7580c2",
  1335 => x"38777a25",
  1336 => x"a138771b",
  1337 => x"70337081",
  1338 => x"ff065858",
  1339 => x"59758a2e",
  1340 => x"98387681",
  1341 => x"ff0651df",
  1342 => x"cb3f8118",
  1343 => x"58797824",
  1344 => x"e13879b0",
  1345 => x"0c8d3d0d",
  1346 => x"048d51df",
  1347 => x"b73f7833",
  1348 => x"7081ff06",
  1349 => x"5257dfac",
  1350 => x"3f811858",
  1351 => x"e0397955",
  1352 => x"7a547d53",
  1353 => x"85528d3d",
  1354 => x"fc0551de",
  1355 => x"943fb008",
  1356 => x"56868b3f",
  1357 => x"7bb0080c",
  1358 => x"75b00c8d",
  1359 => x"3d0d04f6",
  1360 => x"3d0d7d7f",
  1361 => x"80c8bc08",
  1362 => x"705b585a",
  1363 => x"5a7580c1",
  1364 => x"38777925",
  1365 => x"b338dec7",
  1366 => x"3fb00881",
  1367 => x"ff06708d",
  1368 => x"32703070",
  1369 => x"9f2a5151",
  1370 => x"5757768a",
  1371 => x"2e80c338",
  1372 => x"75802ebe",
  1373 => x"38771a56",
  1374 => x"76763476",
  1375 => x"51dec53f",
  1376 => x"81185878",
  1377 => x"7824cf38",
  1378 => x"775675b0",
  1379 => x"0c8c3d0d",
  1380 => x"04785579",
  1381 => x"547c5384",
  1382 => x"528c3dfc",
  1383 => x"0551dda1",
  1384 => x"3fb00856",
  1385 => x"85983f7a",
  1386 => x"b0080c75",
  1387 => x"b00c8c3d",
  1388 => x"0d04771a",
  1389 => x"568a7634",
  1390 => x"8118588d",
  1391 => x"51de853f",
  1392 => x"8a51de80",
  1393 => x"3f7756c2",
  1394 => x"39f93d0d",
  1395 => x"795780c8",
  1396 => x"bc08802e",
  1397 => x"ac387651",
  1398 => x"879e3f7b",
  1399 => x"567a55b0",
  1400 => x"08810554",
  1401 => x"76538252",
  1402 => x"893dfc05",
  1403 => x"51dcd23f",
  1404 => x"b0085784",
  1405 => x"c93f77b0",
  1406 => x"080c76b0",
  1407 => x"0c893d0d",
  1408 => x"0484bb3f",
  1409 => x"850bb008",
  1410 => x"0cff0bb0",
  1411 => x"0c893d0d",
  1412 => x"04fb3d0d",
  1413 => x"80c8bc08",
  1414 => x"70565473",
  1415 => x"883874b0",
  1416 => x"0c873d0d",
  1417 => x"04775383",
  1418 => x"52873dfc",
  1419 => x"0551dc91",
  1420 => x"3fb00854",
  1421 => x"84883f75",
  1422 => x"b0080c73",
  1423 => x"b00c873d",
  1424 => x"0d04ff0b",
  1425 => x"b00c04fb",
  1426 => x"3d0d7755",
  1427 => x"80c8bc08",
  1428 => x"802ea838",
  1429 => x"745186a0",
  1430 => x"3fb00881",
  1431 => x"05547453",
  1432 => x"8752873d",
  1433 => x"fc0551db",
  1434 => x"d83fb008",
  1435 => x"5583cf3f",
  1436 => x"75b0080c",
  1437 => x"74b00c87",
  1438 => x"3d0d0483",
  1439 => x"c13f850b",
  1440 => x"b0080cff",
  1441 => x"0bb00c87",
  1442 => x"3d0d04fa",
  1443 => x"3d0d80c8",
  1444 => x"bc08802e",
  1445 => x"a2387a55",
  1446 => x"79547853",
  1447 => x"8652883d",
  1448 => x"fc0551db",
  1449 => x"9c3fb008",
  1450 => x"5683933f",
  1451 => x"76b0080c",
  1452 => x"75b00c88",
  1453 => x"3d0d0483",
  1454 => x"853f9d0b",
  1455 => x"b0080cff",
  1456 => x"0bb00c88",
  1457 => x"3d0d04fb",
  1458 => x"3d0d7779",
  1459 => x"56568070",
  1460 => x"54547375",
  1461 => x"259f3874",
  1462 => x"101010f8",
  1463 => x"05527216",
  1464 => x"70337074",
  1465 => x"2b760781",
  1466 => x"16f81656",
  1467 => x"56565151",
  1468 => x"747324ea",
  1469 => x"3873b00c",
  1470 => x"873d0d04",
  1471 => x"fc3d0d76",
  1472 => x"785555bc",
  1473 => x"53805273",
  1474 => x"5183de3f",
  1475 => x"84527451",
  1476 => x"ffb53fb0",
  1477 => x"08742384",
  1478 => x"52841551",
  1479 => x"ffa93fb0",
  1480 => x"08821523",
  1481 => x"84528815",
  1482 => x"51ff9c3f",
  1483 => x"b0088415",
  1484 => x"0c84528c",
  1485 => x"1551ff8f",
  1486 => x"3fb00888",
  1487 => x"15238452",
  1488 => x"901551ff",
  1489 => x"823fb008",
  1490 => x"8a152384",
  1491 => x"52941551",
  1492 => x"fef53fb0",
  1493 => x"088c1523",
  1494 => x"84529815",
  1495 => x"51fee83f",
  1496 => x"b0088e15",
  1497 => x"2388529c",
  1498 => x"1551fedb",
  1499 => x"3fb00890",
  1500 => x"150c863d",
  1501 => x"0d04e93d",
  1502 => x"0d6a80c8",
  1503 => x"bc085757",
  1504 => x"75933880",
  1505 => x"c0800b84",
  1506 => x"180c75ac",
  1507 => x"180c75b0",
  1508 => x"0c993d0d",
  1509 => x"04893d70",
  1510 => x"556a5455",
  1511 => x"8a52993d",
  1512 => x"ffbc0551",
  1513 => x"d99b3fb0",
  1514 => x"08775375",
  1515 => x"5256fecc",
  1516 => x"3f818b3f",
  1517 => x"77b0080c",
  1518 => x"75b00c99",
  1519 => x"3d0d04e9",
  1520 => x"3d0d6957",
  1521 => x"80c8bc08",
  1522 => x"802eb538",
  1523 => x"765183a8",
  1524 => x"3f893d70",
  1525 => x"56b00881",
  1526 => x"05557754",
  1527 => x"568f5299",
  1528 => x"3dffbc05",
  1529 => x"51d8da3f",
  1530 => x"b0086b53",
  1531 => x"765257fe",
  1532 => x"8b3f80ca",
  1533 => x"3f77b008",
  1534 => x"0c76b00c",
  1535 => x"993d0d04",
  1536 => x"bd3f850b",
  1537 => x"b0080cff",
  1538 => x"0bb00c99",
  1539 => x"3d0d04fc",
  1540 => x"3d0d8154",
  1541 => x"80c8bc08",
  1542 => x"883873b0",
  1543 => x"0c863d0d",
  1544 => x"04765397",
  1545 => x"b952863d",
  1546 => x"fc0551d8",
  1547 => x"943fb008",
  1548 => x"548c3f74",
  1549 => x"b0080c73",
  1550 => x"b00c863d",
  1551 => x"0d0480c0",
  1552 => x"c808b00c",
  1553 => x"04f73d0d",
  1554 => x"7b80c0c8",
  1555 => x"0882c811",
  1556 => x"085a545a",
  1557 => x"77802e80",
  1558 => x"da388188",
  1559 => x"18841908",
  1560 => x"ff058171",
  1561 => x"2b595559",
  1562 => x"80742480",
  1563 => x"ea388074",
  1564 => x"24b53873",
  1565 => x"822b7811",
  1566 => x"88055656",
  1567 => x"81801908",
  1568 => x"77065372",
  1569 => x"802eb638",
  1570 => x"78167008",
  1571 => x"53537951",
  1572 => x"74085372",
  1573 => x"2dff14fc",
  1574 => x"17fc1779",
  1575 => x"812c5a57",
  1576 => x"57547380",
  1577 => x"25d63877",
  1578 => x"085877ff",
  1579 => x"ad3880c0",
  1580 => x"c80853bc",
  1581 => x"1308a538",
  1582 => x"7951f889",
  1583 => x"3f740853",
  1584 => x"722dff14",
  1585 => x"fc17fc17",
  1586 => x"79812c5a",
  1587 => x"57575473",
  1588 => x"8025ffa8",
  1589 => x"38d13980",
  1590 => x"57ff9339",
  1591 => x"7251bc13",
  1592 => x"0853722d",
  1593 => x"7951f7dd",
  1594 => x"3ffc3d0d",
  1595 => x"76797102",
  1596 => x"8c059f05",
  1597 => x"33575553",
  1598 => x"55837227",
  1599 => x"8a387483",
  1600 => x"06517080",
  1601 => x"2ea238ff",
  1602 => x"125271ff",
  1603 => x"2e933873",
  1604 => x"73708105",
  1605 => x"5534ff12",
  1606 => x"5271ff2e",
  1607 => x"098106ef",
  1608 => x"3874b00c",
  1609 => x"863d0d04",
  1610 => x"7474882b",
  1611 => x"75077071",
  1612 => x"902b0751",
  1613 => x"54518f72",
  1614 => x"27a53872",
  1615 => x"71708405",
  1616 => x"530c7271",
  1617 => x"70840553",
  1618 => x"0c727170",
  1619 => x"8405530c",
  1620 => x"72717084",
  1621 => x"05530cf0",
  1622 => x"1252718f",
  1623 => x"26dd3883",
  1624 => x"72279038",
  1625 => x"72717084",
  1626 => x"05530cfc",
  1627 => x"12527183",
  1628 => x"26f23870",
  1629 => x"53ff9039",
  1630 => x"fd3d0d75",
  1631 => x"70718306",
  1632 => x"53555270",
  1633 => x"b8387170",
  1634 => x"087009f7",
  1635 => x"fbfdff12",
  1636 => x"0670f884",
  1637 => x"82818006",
  1638 => x"51515253",
  1639 => x"709d3884",
  1640 => x"13700870",
  1641 => x"09f7fbfd",
  1642 => x"ff120670",
  1643 => x"f8848281",
  1644 => x"80065151",
  1645 => x"52537080",
  1646 => x"2ee53872",
  1647 => x"52713351",
  1648 => x"70802e8a",
  1649 => x"38811270",
  1650 => x"33525270",
  1651 => x"f8387174",
  1652 => x"31b00c85",
  1653 => x"3d0d04ff",
  1654 => x"3d0d80c7",
  1655 => x"cc0bfc05",
  1656 => x"70085252",
  1657 => x"70ff2e91",
  1658 => x"38702dfc",
  1659 => x"12700852",
  1660 => x"5270ff2e",
  1661 => x"098106f1",
  1662 => x"38833d0d",
  1663 => x"0404d7ad",
  1664 => x"3f040000",
  1665 => x"00ffffff",
  1666 => x"ff00ffff",
  1667 => x"ffff00ff",
  1668 => x"ffffff00",
  1669 => x"00000040",
  1670 => x"44485259",
  1671 => x"53544f4e",
  1672 => x"45205052",
  1673 => x"4f475241",
  1674 => x"4d2c2053",
  1675 => x"4f4d4520",
  1676 => x"53545249",
  1677 => x"4e470000",
  1678 => x"44485259",
  1679 => x"53544f4e",
  1680 => x"45205052",
  1681 => x"4f475241",
  1682 => x"4d2c2031",
  1683 => x"27535420",
  1684 => x"53545249",
  1685 => x"4e470000",
  1686 => x"44687279",
  1687 => x"73746f6e",
  1688 => x"65204265",
  1689 => x"6e63686d",
  1690 => x"61726b2c",
  1691 => x"20566572",
  1692 => x"73696f6e",
  1693 => x"20322e31",
  1694 => x"20284c61",
  1695 => x"6e677561",
  1696 => x"67653a20",
  1697 => x"43290a00",
  1698 => x"50726f67",
  1699 => x"72616d20",
  1700 => x"636f6d70",
  1701 => x"696c6564",
  1702 => x"20776974",
  1703 => x"68202772",
  1704 => x"65676973",
  1705 => x"74657227",
  1706 => x"20617474",
  1707 => x"72696275",
  1708 => x"74650a00",
  1709 => x"45786563",
  1710 => x"7574696f",
  1711 => x"6e207374",
  1712 => x"61727473",
  1713 => x"2c202564",
  1714 => x"2072756e",
  1715 => x"73207468",
  1716 => x"726f7567",
  1717 => x"68204468",
  1718 => x"72797374",
  1719 => x"6f6e650a",
  1720 => x"00000000",
  1721 => x"44485259",
  1722 => x"53544f4e",
  1723 => x"45205052",
  1724 => x"4f475241",
  1725 => x"4d2c2032",
  1726 => x"274e4420",
  1727 => x"53545249",
  1728 => x"4e470000",
  1729 => x"45786563",
  1730 => x"7574696f",
  1731 => x"6e20656e",
  1732 => x"64730a00",
  1733 => x"46696e61",
  1734 => x"6c207661",
  1735 => x"6c756573",
  1736 => x"206f6620",
  1737 => x"74686520",
  1738 => x"76617269",
  1739 => x"61626c65",
  1740 => x"73207573",
  1741 => x"65642069",
  1742 => x"6e207468",
  1743 => x"65206265",
  1744 => x"6e63686d",
  1745 => x"61726b3a",
  1746 => x"0a000000",
  1747 => x"496e745f",
  1748 => x"476c6f62",
  1749 => x"3a202020",
  1750 => x"20202020",
  1751 => x"20202020",
  1752 => x"2025640a",
  1753 => x"00000000",
  1754 => x"20202020",
  1755 => x"20202020",
  1756 => x"73686f75",
  1757 => x"6c642062",
  1758 => x"653a2020",
  1759 => x"2025640a",
  1760 => x"00000000",
  1761 => x"426f6f6c",
  1762 => x"5f476c6f",
  1763 => x"623a2020",
  1764 => x"20202020",
  1765 => x"20202020",
  1766 => x"2025640a",
  1767 => x"00000000",
  1768 => x"43685f31",
  1769 => x"5f476c6f",
  1770 => x"623a2020",
  1771 => x"20202020",
  1772 => x"20202020",
  1773 => x"2025630a",
  1774 => x"00000000",
  1775 => x"20202020",
  1776 => x"20202020",
  1777 => x"73686f75",
  1778 => x"6c642062",
  1779 => x"653a2020",
  1780 => x"2025630a",
  1781 => x"00000000",
  1782 => x"43685f32",
  1783 => x"5f476c6f",
  1784 => x"623a2020",
  1785 => x"20202020",
  1786 => x"20202020",
  1787 => x"2025630a",
  1788 => x"00000000",
  1789 => x"4172725f",
  1790 => x"315f476c",
  1791 => x"6f625b38",
  1792 => x"5d3a2020",
  1793 => x"20202020",
  1794 => x"2025640a",
  1795 => x"00000000",
  1796 => x"4172725f",
  1797 => x"325f476c",
  1798 => x"6f625b38",
  1799 => x"5d5b375d",
  1800 => x"3a202020",
  1801 => x"2025640a",
  1802 => x"00000000",
  1803 => x"20202020",
  1804 => x"20202020",
  1805 => x"73686f75",
  1806 => x"6c642062",
  1807 => x"653a2020",
  1808 => x"204e756d",
  1809 => x"6265725f",
  1810 => x"4f665f52",
  1811 => x"756e7320",
  1812 => x"2b203130",
  1813 => x"0a000000",
  1814 => x"5074725f",
  1815 => x"476c6f62",
  1816 => x"2d3e0a00",
  1817 => x"20205074",
  1818 => x"725f436f",
  1819 => x"6d703a20",
  1820 => x"20202020",
  1821 => x"20202020",
  1822 => x"2025640a",
  1823 => x"00000000",
  1824 => x"20202020",
  1825 => x"20202020",
  1826 => x"73686f75",
  1827 => x"6c642062",
  1828 => x"653a2020",
  1829 => x"2028696d",
  1830 => x"706c656d",
  1831 => x"656e7461",
  1832 => x"74696f6e",
  1833 => x"2d646570",
  1834 => x"656e6465",
  1835 => x"6e74290a",
  1836 => x"00000000",
  1837 => x"20204469",
  1838 => x"7363723a",
  1839 => x"20202020",
  1840 => x"20202020",
  1841 => x"20202020",
  1842 => x"2025640a",
  1843 => x"00000000",
  1844 => x"2020456e",
  1845 => x"756d5f43",
  1846 => x"6f6d703a",
  1847 => x"20202020",
  1848 => x"20202020",
  1849 => x"2025640a",
  1850 => x"00000000",
  1851 => x"2020496e",
  1852 => x"745f436f",
  1853 => x"6d703a20",
  1854 => x"20202020",
  1855 => x"20202020",
  1856 => x"2025640a",
  1857 => x"00000000",
  1858 => x"20205374",
  1859 => x"725f436f",
  1860 => x"6d703a20",
  1861 => x"20202020",
  1862 => x"20202020",
  1863 => x"2025730a",
  1864 => x"00000000",
  1865 => x"20202020",
  1866 => x"20202020",
  1867 => x"73686f75",
  1868 => x"6c642062",
  1869 => x"653a2020",
  1870 => x"20444852",
  1871 => x"5953544f",
  1872 => x"4e452050",
  1873 => x"524f4752",
  1874 => x"414d2c20",
  1875 => x"534f4d45",
  1876 => x"20535452",
  1877 => x"494e470a",
  1878 => x"00000000",
  1879 => x"4e657874",
  1880 => x"5f507472",
  1881 => x"5f476c6f",
  1882 => x"622d3e0a",
  1883 => x"00000000",
  1884 => x"20202020",
  1885 => x"20202020",
  1886 => x"73686f75",
  1887 => x"6c642062",
  1888 => x"653a2020",
  1889 => x"2028696d",
  1890 => x"706c656d",
  1891 => x"656e7461",
  1892 => x"74696f6e",
  1893 => x"2d646570",
  1894 => x"656e6465",
  1895 => x"6e74292c",
  1896 => x"2073616d",
  1897 => x"65206173",
  1898 => x"2061626f",
  1899 => x"76650a00",
  1900 => x"496e745f",
  1901 => x"315f4c6f",
  1902 => x"633a2020",
  1903 => x"20202020",
  1904 => x"20202020",
  1905 => x"2025640a",
  1906 => x"00000000",
  1907 => x"496e745f",
  1908 => x"325f4c6f",
  1909 => x"633a2020",
  1910 => x"20202020",
  1911 => x"20202020",
  1912 => x"2025640a",
  1913 => x"00000000",
  1914 => x"496e745f",
  1915 => x"335f4c6f",
  1916 => x"633a2020",
  1917 => x"20202020",
  1918 => x"20202020",
  1919 => x"2025640a",
  1920 => x"00000000",
  1921 => x"456e756d",
  1922 => x"5f4c6f63",
  1923 => x"3a202020",
  1924 => x"20202020",
  1925 => x"20202020",
  1926 => x"2025640a",
  1927 => x"00000000",
  1928 => x"5374725f",
  1929 => x"315f4c6f",
  1930 => x"633a2020",
  1931 => x"20202020",
  1932 => x"20202020",
  1933 => x"2025730a",
  1934 => x"00000000",
  1935 => x"20202020",
  1936 => x"20202020",
  1937 => x"73686f75",
  1938 => x"6c642062",
  1939 => x"653a2020",
  1940 => x"20444852",
  1941 => x"5953544f",
  1942 => x"4e452050",
  1943 => x"524f4752",
  1944 => x"414d2c20",
  1945 => x"31275354",
  1946 => x"20535452",
  1947 => x"494e470a",
  1948 => x"00000000",
  1949 => x"5374725f",
  1950 => x"325f4c6f",
  1951 => x"633a2020",
  1952 => x"20202020",
  1953 => x"20202020",
  1954 => x"2025730a",
  1955 => x"00000000",
  1956 => x"20202020",
  1957 => x"20202020",
  1958 => x"73686f75",
  1959 => x"6c642062",
  1960 => x"653a2020",
  1961 => x"20444852",
  1962 => x"5953544f",
  1963 => x"4e452050",
  1964 => x"524f4752",
  1965 => x"414d2c20",
  1966 => x"32274e44",
  1967 => x"20535452",
  1968 => x"494e470a",
  1969 => x"00000000",
  1970 => x"55736572",
  1971 => x"2074696d",
  1972 => x"653a2025",
  1973 => x"640a0000",
  1974 => x"4d696372",
  1975 => x"6f736563",
  1976 => x"6f6e6473",
  1977 => x"20666f72",
  1978 => x"206f6e65",
  1979 => x"2072756e",
  1980 => x"20746872",
  1981 => x"6f756768",
  1982 => x"20446872",
  1983 => x"7973746f",
  1984 => x"6e653a20",
  1985 => x"00000000",
  1986 => x"2564200a",
  1987 => x"00000000",
  1988 => x"44687279",
  1989 => x"73746f6e",
  1990 => x"65732070",
  1991 => x"65722053",
  1992 => x"65636f6e",
  1993 => x"643a2020",
  1994 => x"20202020",
  1995 => x"20202020",
  1996 => x"20202020",
  1997 => x"20202020",
  1998 => x"20202020",
  1999 => x"00000000",
  2000 => x"56415820",
  2001 => x"4d495053",
  2002 => x"20726174",
  2003 => x"696e6720",
  2004 => x"2a203130",
  2005 => x"3030203d",
  2006 => x"20256420",
  2007 => x"0a000000",
  2008 => x"50726f67",
  2009 => x"72616d20",
  2010 => x"636f6d70",
  2011 => x"696c6564",
  2012 => x"20776974",
  2013 => x"686f7574",
  2014 => x"20277265",
  2015 => x"67697374",
  2016 => x"65722720",
  2017 => x"61747472",
  2018 => x"69627574",
  2019 => x"650a0000",
  2020 => x"4d656173",
  2021 => x"75726564",
  2022 => x"2074696d",
  2023 => x"6520746f",
  2024 => x"6f20736d",
  2025 => x"616c6c20",
  2026 => x"746f206f",
  2027 => x"62746169",
  2028 => x"6e206d65",
  2029 => x"616e696e",
  2030 => x"6766756c",
  2031 => x"20726573",
  2032 => x"756c7473",
  2033 => x"0a000000",
  2034 => x"506c6561",
  2035 => x"73652069",
  2036 => x"6e637265",
  2037 => x"61736520",
  2038 => x"6e756d62",
  2039 => x"6572206f",
  2040 => x"66207275",
  2041 => x"6e730a00",
  2042 => x"44485259",
  2043 => x"53544f4e",
  2044 => x"45205052",
  2045 => x"4f475241",
  2046 => x"4d2c2033",
  2047 => x"27524420",
  2048 => x"53545249",
  2049 => x"4e470000",
  2050 => x"30313233",
  2051 => x"34353637",
  2052 => x"38394142",
  2053 => x"43444546",
  2054 => x"00000000",
  2055 => x"64756d6d",
  2056 => x"792e6578",
  2057 => x"65000000",
  2058 => x"43000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"000023d4",
  2063 => x"000061a8",
  2064 => x"00000000",
  2065 => x"0000201c",
  2066 => x"0000204c",
  2067 => x"00000000",
  2068 => x"000022b4",
  2069 => x"00002310",
  2070 => x"0000236c",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00002028",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000001",
  2110 => x"330eabcd",
  2111 => x"1234e66d",
  2112 => x"deec0005",
  2113 => x"000b0000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"00000000",
  2209 => x"00000000",
  2210 => x"00000000",
  2211 => x"00000000",
  2212 => x"00000000",
  2213 => x"00000000",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"00000000",
  2217 => x"00000000",
  2218 => x"00000000",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000000",
  2244 => x"00000000",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"00000000",
  2262 => x"00000000",
  2263 => x"00000000",
  2264 => x"00000000",
  2265 => x"00000000",
  2266 => x"00000000",
  2267 => x"00000000",
  2268 => x"00000000",
  2269 => x"00000000",
  2270 => x"00000000",
  2271 => x"00000000",
  2272 => x"00000000",
  2273 => x"00000000",
  2274 => x"00000000",
  2275 => x"00000000",
  2276 => x"00000000",
  2277 => x"00000000",
  2278 => x"00000000",
  2279 => x"00000000",
  2280 => x"00000000",
  2281 => x"00000000",
  2282 => x"00000000",
  2283 => x"00000000",
  2284 => x"00000000",
  2285 => x"00000000",
  2286 => x"00000000",
  2287 => x"00000000",
  2288 => x"00000000",
  2289 => x"00000000",
  2290 => x"ffffffff",
  2291 => x"00000000",
  2292 => x"ffffffff",
  2293 => x"00000000",
  2294 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;


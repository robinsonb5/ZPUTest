-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity sdbootstrap_rom is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end sdbootstrap_rom;

architecture arch of sdbootstrap_rom is
begin

type ram_type is array(natural range 0 to ((2**(maxAddrBitStackBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(

     0 => x"a08080f4",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"9cb87383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02ec050d",
    30 => x"88bd0bff",
    31 => x"880c800b",
    32 => x"870a0cf8",
    33 => x"0883fff0",
    34 => x"900cfc08",
    35 => x"83fff094",
    36 => x"0c84eacd",
    37 => x"a8800b83",
    38 => x"fff0980c",
    39 => x"a0808790",
    40 => x"2d83ffe0",
    41 => x"8008902b",
    42 => x"70902c51",
    43 => x"5372802e",
    44 => x"81d138a0",
    45 => x"808f822d",
    46 => x"83ffe090",
    47 => x"5283fff0",
    48 => x"9051a080",
    49 => x"9a932d83",
    50 => x"ffe08008",
    51 => x"802e81b3",
    52 => x"3883ffe0",
    53 => x"90548055",
    54 => x"73708105",
    55 => x"55a08080",
    56 => x"b42d5372",
    57 => x"a02e80de",
    58 => x"3872a32e",
    59 => x"80fd3872",
    60 => x"80c72e09",
    61 => x"81068b38",
    62 => x"a0808088",
    63 => x"2da08082",
    64 => x"a204728a",
    65 => x"2e098106",
    66 => x"8b38a080",
    67 => x"80902da0",
    68 => x"8082a204",
    69 => x"7280cc2e",
    70 => x"09810686",
    71 => x"3883ffe0",
    72 => x"90547281",
    73 => x"df06f005",
    74 => x"7081ff06",
    75 => x"5153b873",
    76 => x"278938ef",
    77 => x"137081ff",
    78 => x"06515374",
    79 => x"842b7307",
    80 => x"55a08081",
    81 => x"d80472a3",
    82 => x"2ea13873",
    83 => x"70810555",
    84 => x"a08080b4",
    85 => x"2d5372a0",
    86 => x"2ef138ff",
    87 => x"14755370",
    88 => x"5254a080",
    89 => x"9a932d74",
    90 => x"870a0c73",
    91 => x"70810555",
    92 => x"a08080b4",
    93 => x"2d53728a",
    94 => x"2e098106",
    95 => x"ee38a080",
    96 => x"81d60480",
    97 => x"0b83ffe0",
    98 => x"800c0294",
    99 => x"050d0402",
   100 => x"f4050d74",
   101 => x"767181ff",
   102 => x"06c80c53",
   103 => x"5383fff0",
   104 => x"9c088538",
   105 => x"71892b52",
   106 => x"71982ac8",
   107 => x"0c71902a",
   108 => x"7081ff06",
   109 => x"c80c5171",
   110 => x"882a7081",
   111 => x"ff06c80c",
   112 => x"517181ff",
   113 => x"06c80c72",
   114 => x"902a7081",
   115 => x"ff06c80c",
   116 => x"51c80870",
   117 => x"81ff0651",
   118 => x"5182b8bf",
   119 => x"527081ff",
   120 => x"2e098106",
   121 => x"943881ff",
   122 => x"0bc80cc8",
   123 => x"087081ff",
   124 => x"06ff1454",
   125 => x"515171e5",
   126 => x"387083ff",
   127 => x"e0800c02",
   128 => x"8c050d04",
   129 => x"02fc050d",
   130 => x"81c75181",
   131 => x"ff0bc80c",
   132 => x"ff115170",
   133 => x"8025f438",
   134 => x"0284050d",
   135 => x"0402ec05",
   136 => x"0da08084",
   137 => x"842d819c",
   138 => x"9f558052",
   139 => x"87fc80f7",
   140 => x"51a08083",
   141 => x"8f2d83ff",
   142 => x"e0800890",
   143 => x"2b70902c",
   144 => x"70565153",
   145 => x"72812e09",
   146 => x"8106b338",
   147 => x"81ff0bc8",
   148 => x"0c820a52",
   149 => x"849c80e9",
   150 => x"51a08083",
   151 => x"8f2d83ff",
   152 => x"e0800890",
   153 => x"2b70902c",
   154 => x"5153728d",
   155 => x"3881ff0b",
   156 => x"c80c7353",
   157 => x"a0808587",
   158 => x"04a08084",
   159 => x"842dff15",
   160 => x"5574ffa6",
   161 => x"38745372",
   162 => x"83ffe080",
   163 => x"0c029405",
   164 => x"0d0402f0",
   165 => x"050d81ff",
   166 => x"0bc80c93",
   167 => x"54805287",
   168 => x"fc80c151",
   169 => x"a080838f",
   170 => x"2d83ffe0",
   171 => x"8008902b",
   172 => x"70902c51",
   173 => x"53728d38",
   174 => x"81ff0bc8",
   175 => x"0c8153a0",
   176 => x"8085d104",
   177 => x"a0808484",
   178 => x"2dff1454",
   179 => x"73cf3873",
   180 => x"537283ff",
   181 => x"e0800c02",
   182 => x"90050d04",
   183 => x"02f0050d",
   184 => x"a0808484",
   185 => x"2d83aa52",
   186 => x"849c80c8",
   187 => x"51a08083",
   188 => x"8f2d83ff",
   189 => x"e0800881",
   190 => x"2e098106",
   191 => x"9038cc08",
   192 => x"7083ffff",
   193 => x"06515372",
   194 => x"83aa2e99",
   195 => x"38a08085",
   196 => x"922da080",
   197 => x"869e0481",
   198 => x"54a08087",
   199 => x"85048054",
   200 => x"a0808785",
   201 => x"0481ff0b",
   202 => x"c80cb154",
   203 => x"a080849d",
   204 => x"2d83ffe0",
   205 => x"8008902b",
   206 => x"70902c51",
   207 => x"5372802e",
   208 => x"b7388052",
   209 => x"87fc80fa",
   210 => x"51a08083",
   211 => x"8f2d83ff",
   212 => x"e08008a4",
   213 => x"3881ff0b",
   214 => x"c80cc808",
   215 => x"cc087186",
   216 => x"2a708106",
   217 => x"83ffe080",
   218 => x"08535152",
   219 => x"55537280",
   220 => x"2e9338a0",
   221 => x"80869704",
   222 => x"73822eff",
   223 => x"a138ff14",
   224 => x"5473ffa8",
   225 => x"387383ff",
   226 => x"e0800c02",
   227 => x"90050d04",
   228 => x"02f4050d",
   229 => x"810b83ff",
   230 => x"f09c0cc4",
   231 => x"08708f2a",
   232 => x"70810651",
   233 => x"515372f3",
   234 => x"3872c40c",
   235 => x"a0808484",
   236 => x"2dc40870",
   237 => x"8f2a7081",
   238 => x"06515153",
   239 => x"72f33881",
   240 => x"0bc40c87",
   241 => x"53805284",
   242 => x"d480c051",
   243 => x"a080838f",
   244 => x"2d83ffe0",
   245 => x"8008812e",
   246 => x"96387282",
   247 => x"2e098106",
   248 => x"88388053",
   249 => x"a08088ad",
   250 => x"04ff1353",
   251 => x"72d738a0",
   252 => x"8085dc2d",
   253 => x"83ffe080",
   254 => x"08902b70",
   255 => x"902c83ff",
   256 => x"f09c0c53",
   257 => x"815287fc",
   258 => x"80d051a0",
   259 => x"80838f2d",
   260 => x"81ff0bc8",
   261 => x"0cc40870",
   262 => x"8f2a7081",
   263 => x"06515153",
   264 => x"72f33872",
   265 => x"c40c81ff",
   266 => x"0bc80c81",
   267 => x"537283ff",
   268 => x"e0800c02",
   269 => x"8c050d04",
   270 => x"800b83ff",
   271 => x"e0800c04",
   272 => x"02e8050d",
   273 => x"78558056",
   274 => x"c408708f",
   275 => x"2a708106",
   276 => x"51515372",
   277 => x"f3388281",
   278 => x"0bc40c81",
   279 => x"ff0bc80c",
   280 => x"775287fc",
   281 => x"80d151a0",
   282 => x"80838f2d",
   283 => x"83ffe080",
   284 => x"0880d238",
   285 => x"80dbc6df",
   286 => x"5481ff0b",
   287 => x"c80cc808",
   288 => x"7081ff06",
   289 => x"51537281",
   290 => x"fe2e0981",
   291 => x"069b3880",
   292 => x"ff54cc08",
   293 => x"75708405",
   294 => x"570cff14",
   295 => x"54738025",
   296 => x"f1388156",
   297 => x"a08089af",
   298 => x"04ff1454",
   299 => x"73cb3881",
   300 => x"ff0bc80c",
   301 => x"c408708f",
   302 => x"2a708106",
   303 => x"51515372",
   304 => x"f33872c4",
   305 => x"0c7583ff",
   306 => x"e0800c02",
   307 => x"98050d04",
   308 => x"02e0050d",
   309 => x"795683ff",
   310 => x"fe800b83",
   311 => x"fff0bc0c",
   312 => x"83fffe80",
   313 => x"528051a0",
   314 => x"8088c02d",
   315 => x"83ffe080",
   316 => x"08902b70",
   317 => x"902c7056",
   318 => x"51537280",
   319 => x"2e839c38",
   320 => x"83fff0bc",
   321 => x"0883fe11",
   322 => x"a08080b4",
   323 => x"2d545572",
   324 => x"80d52e09",
   325 => x"810681f8",
   326 => x"3883ff15",
   327 => x"a08080b4",
   328 => x"2d537281",
   329 => x"aa2e0981",
   330 => x"0681e538",
   331 => x"7580f038",
   332 => x"83be158b",
   333 => x"11a08080",
   334 => x"b42d8a12",
   335 => x"a08080b4",
   336 => x"2d71982b",
   337 => x"71902b07",
   338 => x"8914a080",
   339 => x"80b42d70",
   340 => x"882b7207",
   341 => x"8816a080",
   342 => x"80b42d71",
   343 => x"077083ff",
   344 => x"f0c00c7b",
   345 => x"59575253",
   346 => x"575a5853",
   347 => x"a08088c0",
   348 => x"2d83fff0",
   349 => x"bc0883fe",
   350 => x"11a08080",
   351 => x"b42d5454",
   352 => x"7280d52e",
   353 => x"09810690",
   354 => x"3883ff14",
   355 => x"a08080b4",
   356 => x"2d537281",
   357 => x"aa2e8838",
   358 => x"7554a080",
   359 => x"8d9b0480",
   360 => x"0b83fff0",
   361 => x"ac0c83ff",
   362 => x"f0bc08b6",
   363 => x"11545572",
   364 => x"0884b285",
   365 => x"a8b12e09",
   366 => x"8106ab38",
   367 => x"84130883",
   368 => x"9180c0a0",
   369 => x"2e098106",
   370 => x"88388c0b",
   371 => x"83fff0ac",
   372 => x"0c841308",
   373 => x"83b180c0",
   374 => x"a02e0981",
   375 => x"06883890",
   376 => x"0b83fff0",
   377 => x"ac0c83ff",
   378 => x"f0ac0870",
   379 => x"55567580",
   380 => x"2e81a838",
   381 => x"88158311",
   382 => x"a08080b4",
   383 => x"2d585376",
   384 => x"8f388413",
   385 => x"0883fe80",
   386 => x"06537284",
   387 => x"802e8838",
   388 => x"8054a080",
   389 => x"8d9b048f",
   390 => x"15a08080",
   391 => x"b42d8e16",
   392 => x"a08080b4",
   393 => x"2d71882b",
   394 => x"0783fff0",
   395 => x"a8080570",
   396 => x"83fff0a8",
   397 => x"0c555875",
   398 => x"8c2e8a38",
   399 => x"75902e09",
   400 => x"810680d7",
   401 => x"387683ff",
   402 => x"f0b00c73",
   403 => x"83fff0b4",
   404 => x"0c9115a0",
   405 => x"8080b42d",
   406 => x"9016a080",
   407 => x"80b42d71",
   408 => x"882b078a",
   409 => x"17a08080",
   410 => x"b42dff05",
   411 => x"55575772",
   412 => x"802e9038",
   413 => x"7514ff14",
   414 => x"545472f8",
   415 => x"387383ff",
   416 => x"f0b40c8c",
   417 => x"15a08080",
   418 => x"b42d8b16",
   419 => x"a08080b4",
   420 => x"2d71882b",
   421 => x"0783fff0",
   422 => x"b80c5873",
   423 => x"83ffe080",
   424 => x"0c02a005",
   425 => x"0d0402fc",
   426 => x"050d7083",
   427 => x"ffe0800c",
   428 => x"0284050d",
   429 => x"0402fc05",
   430 => x"0d7083ff",
   431 => x"e0800c02",
   432 => x"84050d04",
   433 => x"02fc050d",
   434 => x"7083ffe0",
   435 => x"800c0284",
   436 => x"050d0402",
   437 => x"f8050d81",
   438 => x"51a08089",
   439 => x"d02d83ff",
   440 => x"e080089b",
   441 => x"3883ffe0",
   442 => x"800851a0",
   443 => x"8089d02d",
   444 => x"83ffe080",
   445 => x"085283ff",
   446 => x"e0800880",
   447 => x"2eb138a0",
   448 => x"808da62d",
   449 => x"83ffe080",
   450 => x"08802ea1",
   451 => x"387351a0",
   452 => x"808db52d",
   453 => x"83ffe080",
   454 => x"08802e91",
   455 => x"387451a0",
   456 => x"808dc42d",
   457 => x"815283ff",
   458 => x"e0800883",
   459 => x"38805271",
   460 => x"83ffe080",
   461 => x"0c028805",
   462 => x"0d0402e8",
   463 => x"050d7779",
   464 => x"7b585555",
   465 => x"80537276",
   466 => x"25ab3874",
   467 => x"70810556",
   468 => x"a08080b4",
   469 => x"2d747081",
   470 => x"0556a080",
   471 => x"80b42d52",
   472 => x"5271712e",
   473 => x"88388151",
   474 => x"a0808ef7",
   475 => x"04811353",
   476 => x"a0808ec6",
   477 => x"04805170",
   478 => x"83ffe080",
   479 => x"0c029805",
   480 => x"0d0402d8",
   481 => x"050dff0b",
   482 => x"83fff4e4",
   483 => x"0c800b83",
   484 => x"fff4f80c",
   485 => x"83fff0d0",
   486 => x"528051a0",
   487 => x"8088c02d",
   488 => x"83ffe080",
   489 => x"08902b70",
   490 => x"902c7057",
   491 => x"51547380",
   492 => x"2e86d738",
   493 => x"8056810b",
   494 => x"83fff0c4",
   495 => x"0c8853a0",
   496 => x"809cc852",
   497 => x"83fff186",
   498 => x"51a0808e",
   499 => x"ba2d83ff",
   500 => x"e0800876",
   501 => x"2e098106",
   502 => x"8b3883ff",
   503 => x"e0800883",
   504 => x"fff0c40c",
   505 => x"8853a080",
   506 => x"9cd45283",
   507 => x"fff1a251",
   508 => x"a0808eba",
   509 => x"2d83ffe0",
   510 => x"80088b38",
   511 => x"83ffe080",
   512 => x"0883fff0",
   513 => x"c40c83ff",
   514 => x"f0c40880",
   515 => x"2e81a038",
   516 => x"83fff496",
   517 => x"0ba08080",
   518 => x"b42d83ff",
   519 => x"f4970ba0",
   520 => x"8080b42d",
   521 => x"71982b71",
   522 => x"902b0783",
   523 => x"fff4980b",
   524 => x"a08080b4",
   525 => x"2d70882b",
   526 => x"720783ff",
   527 => x"f4990ba0",
   528 => x"8080b42d",
   529 => x"710783ff",
   530 => x"f4ce0ba0",
   531 => x"8080b42d",
   532 => x"83fff4cf",
   533 => x"0ba08080",
   534 => x"b42d7188",
   535 => x"2b07535f",
   536 => x"54525a56",
   537 => x"57557381",
   538 => x"abaa2e09",
   539 => x"81069338",
   540 => x"7551a080",
   541 => x"9bc92d83",
   542 => x"ffe08008",
   543 => x"56a08091",
   544 => x"8f048055",
   545 => x"7382d4d5",
   546 => x"2e098106",
   547 => x"84fc3883",
   548 => x"fff0d052",
   549 => x"7551a080",
   550 => x"88c02d83",
   551 => x"ffe08008",
   552 => x"902b7090",
   553 => x"2c705751",
   554 => x"5473802e",
   555 => x"84dc3888",
   556 => x"53a0809c",
   557 => x"d45283ff",
   558 => x"f1a251a0",
   559 => x"808eba2d",
   560 => x"83ffe080",
   561 => x"088d3881",
   562 => x"0b83fff4",
   563 => x"f80ca080",
   564 => x"91f30488",
   565 => x"53a0809c",
   566 => x"c85283ff",
   567 => x"f18651a0",
   568 => x"808eba2d",
   569 => x"805583ff",
   570 => x"e0800875",
   571 => x"2e098106",
   572 => x"84983883",
   573 => x"fff4ce0b",
   574 => x"a08080b4",
   575 => x"2d547380",
   576 => x"d52e0981",
   577 => x"0680db38",
   578 => x"83fff4cf",
   579 => x"0ba08080",
   580 => x"b42d5473",
   581 => x"81aa2e09",
   582 => x"810680c6",
   583 => x"38800b83",
   584 => x"fff0d00b",
   585 => x"a08080b4",
   586 => x"2d565474",
   587 => x"81e92e83",
   588 => x"38815474",
   589 => x"81eb2e8c",
   590 => x"38805573",
   591 => x"752e0981",
   592 => x"0683c738",
   593 => x"83fff0db",
   594 => x"0ba08080",
   595 => x"b42d5574",
   596 => x"913883ff",
   597 => x"f0dc0ba0",
   598 => x"8080b42d",
   599 => x"5473822e",
   600 => x"88388055",
   601 => x"a080968a",
   602 => x"0483fff0",
   603 => x"dd0ba080",
   604 => x"80b42d70",
   605 => x"83fff580",
   606 => x"0cff0583",
   607 => x"fff4f40c",
   608 => x"83fff0de",
   609 => x"0ba08080",
   610 => x"b42d83ff",
   611 => x"f0df0ba0",
   612 => x"8080b42d",
   613 => x"58760577",
   614 => x"82802905",
   615 => x"7083fff4",
   616 => x"e80c83ff",
   617 => x"f0e00ba0",
   618 => x"8080b42d",
   619 => x"7083fff4",
   620 => x"e00c83ff",
   621 => x"f4f80859",
   622 => x"57587680",
   623 => x"2e81df38",
   624 => x"8853a080",
   625 => x"9cd45283",
   626 => x"fff1a251",
   627 => x"a0808eba",
   628 => x"2d83ffe0",
   629 => x"800882b2",
   630 => x"3883fff5",
   631 => x"80087084",
   632 => x"2b83fff4",
   633 => x"d00c7083",
   634 => x"fff4fc0c",
   635 => x"83fff0f5",
   636 => x"0ba08080",
   637 => x"b42d83ff",
   638 => x"f0f40ba0",
   639 => x"8080b42d",
   640 => x"71828029",
   641 => x"0583fff0",
   642 => x"f60ba080",
   643 => x"80b42d70",
   644 => x"84808029",
   645 => x"1283fff0",
   646 => x"f70ba080",
   647 => x"80b42d70",
   648 => x"81800a29",
   649 => x"127083ff",
   650 => x"f0c80c83",
   651 => x"fff4e008",
   652 => x"712983ff",
   653 => x"f4e80805",
   654 => x"7083fff5",
   655 => x"880c83ff",
   656 => x"f0fd0ba0",
   657 => x"8080b42d",
   658 => x"83fff0fc",
   659 => x"0ba08080",
   660 => x"b42d7182",
   661 => x"80290583",
   662 => x"fff0fe0b",
   663 => x"a08080b4",
   664 => x"2d708480",
   665 => x"80291283",
   666 => x"fff0ff0b",
   667 => x"a08080b4",
   668 => x"2d70982b",
   669 => x"81f00a06",
   670 => x"72057083",
   671 => x"fff0cc0c",
   672 => x"fe117e29",
   673 => x"770583ff",
   674 => x"f4f00c52",
   675 => x"59524354",
   676 => x"5e515259",
   677 => x"525d5759",
   678 => x"57a08096",
   679 => x"880483ff",
   680 => x"f0e20ba0",
   681 => x"8080b42d",
   682 => x"83fff0e1",
   683 => x"0ba08080",
   684 => x"b42d7182",
   685 => x"80290570",
   686 => x"83fff4d0",
   687 => x"0c70a029",
   688 => x"83ff0570",
   689 => x"892a7083",
   690 => x"fff4fc0c",
   691 => x"83fff0e7",
   692 => x"0ba08080",
   693 => x"b42d83ff",
   694 => x"f0e60ba0",
   695 => x"8080b42d",
   696 => x"71828029",
   697 => x"057083ff",
   698 => x"f0c80c7b",
   699 => x"71291e70",
   700 => x"83fff4f0",
   701 => x"0c7d83ff",
   702 => x"f0cc0c73",
   703 => x"0583fff5",
   704 => x"880c555e",
   705 => x"51515555",
   706 => x"81557483",
   707 => x"ffe0800c",
   708 => x"02a8050d",
   709 => x"0402e805",
   710 => x"0d777087",
   711 => x"2c7180ff",
   712 => x"06565653",
   713 => x"83fff4f8",
   714 => x"088a3872",
   715 => x"882c7381",
   716 => x"ff065555",
   717 => x"7483fff4",
   718 => x"e4082eac",
   719 => x"3883fff0",
   720 => x"d05283ff",
   721 => x"f4e80815",
   722 => x"51a08088",
   723 => x"c02d83ff",
   724 => x"e0800890",
   725 => x"2b70902c",
   726 => x"70585153",
   727 => x"72802e80",
   728 => x"cb387483",
   729 => x"fff4e40c",
   730 => x"83fff4f8",
   731 => x"08802ea0",
   732 => x"38738429",
   733 => x"83fff0d0",
   734 => x"05700852",
   735 => x"53a0809b",
   736 => x"c92d83ff",
   737 => x"e08008f0",
   738 => x"0a0654a0",
   739 => x"8097aa04",
   740 => x"731083ff",
   741 => x"f0d00570",
   742 => x"a080809f",
   743 => x"2d5253a0",
   744 => x"809bfb2d",
   745 => x"83ffe080",
   746 => x"08547356",
   747 => x"7583ffe0",
   748 => x"800c0298",
   749 => x"050d0402",
   750 => x"cc050d7e",
   751 => x"605e5b80",
   752 => x"56ff0b83",
   753 => x"fff4e40c",
   754 => x"83fff0cc",
   755 => x"0883fff4",
   756 => x"f008565a",
   757 => x"83fff4f8",
   758 => x"08762e8e",
   759 => x"3883fff5",
   760 => x"8008842b",
   761 => x"58a08097",
   762 => x"f20483ff",
   763 => x"f4fc0884",
   764 => x"2b588059",
   765 => x"78782781",
   766 => x"c938788f",
   767 => x"06a01757",
   768 => x"54739538",
   769 => x"83fff0d0",
   770 => x"52745181",
   771 => x"1555a080",
   772 => x"88c02d83",
   773 => x"fff0d056",
   774 => x"8076a080",
   775 => x"80b42d55",
   776 => x"5773772e",
   777 => x"83388157",
   778 => x"7381e52e",
   779 => x"818c3881",
   780 => x"70780655",
   781 => x"5c73802e",
   782 => x"8180388b",
   783 => x"16a08080",
   784 => x"b42d9806",
   785 => x"577680f2",
   786 => x"388b537c",
   787 => x"527551a0",
   788 => x"808eba2d",
   789 => x"83ffe080",
   790 => x"0880df38",
   791 => x"9c160851",
   792 => x"a0809bc9",
   793 => x"2d83ffe0",
   794 => x"8008841c",
   795 => x"0c9a16a0",
   796 => x"80809f2d",
   797 => x"51a0809b",
   798 => x"fb2d83ff",
   799 => x"e0800883",
   800 => x"ffe08008",
   801 => x"555583ff",
   802 => x"f4f80880",
   803 => x"2e9e3894",
   804 => x"16a08080",
   805 => x"9f2d51a0",
   806 => x"809bfb2d",
   807 => x"83ffe080",
   808 => x"08902b83",
   809 => x"fff00a06",
   810 => x"70165154",
   811 => x"73881c0c",
   812 => x"767b0c7b",
   813 => x"54a0809a",
   814 => x"88048119",
   815 => x"59a08097",
   816 => x"f40483ff",
   817 => x"f4f80880",
   818 => x"2ebc3879",
   819 => x"51a08096",
   820 => x"952d83ff",
   821 => x"e0800883",
   822 => x"ffe08008",
   823 => x"80ffffff",
   824 => x"f806555a",
   825 => x"7380ffff",
   826 => x"fff82e9a",
   827 => x"3883ffe0",
   828 => x"8008fe05",
   829 => x"83fff580",
   830 => x"082983ff",
   831 => x"f5880805",
   832 => x"55a08097",
   833 => x"f2048054",
   834 => x"7383ffe0",
   835 => x"800c02b4",
   836 => x"050d0402",
   837 => x"e4050d79",
   838 => x"795383ff",
   839 => x"f4d45255",
   840 => x"a08097b7",
   841 => x"2d83ffe0",
   842 => x"800881ff",
   843 => x"06705553",
   844 => x"72802e81",
   845 => x"893883ff",
   846 => x"f4d80883",
   847 => x"ff05892a",
   848 => x"57807055",
   849 => x"56757725",
   850 => x"80f23883",
   851 => x"fff4dc08",
   852 => x"fe0583ff",
   853 => x"f5800829",
   854 => x"83fff588",
   855 => x"08117583",
   856 => x"fff4f408",
   857 => x"06057654",
   858 => x"5253a080",
   859 => x"88c02d83",
   860 => x"ffe08008",
   861 => x"902b7090",
   862 => x"2c515372",
   863 => x"802eb638",
   864 => x"81147083",
   865 => x"fff4f408",
   866 => x"06545472",
   867 => x"963883ff",
   868 => x"f4dc0851",
   869 => x"a0809695",
   870 => x"2d83ffe0",
   871 => x"800883ff",
   872 => x"f4dc0c84",
   873 => x"80158117",
   874 => x"57557676",
   875 => x"24ff9c38",
   876 => x"a0809bbc",
   877 => x"047254a0",
   878 => x"809bbe04",
   879 => x"81547383",
   880 => x"ffe0800c",
   881 => x"029c050d",
   882 => x"0402f405",
   883 => x"0d747088",
   884 => x"2a83fe80",
   885 => x"06707298",
   886 => x"2a077288",
   887 => x"2b87fc80",
   888 => x"80067398",
   889 => x"2b81f00a",
   890 => x"06717307",
   891 => x"0783ffe0",
   892 => x"800c5651",
   893 => x"5351028c",
   894 => x"050d0402",
   895 => x"f4050d02",
   896 => x"9205a080",
   897 => x"809f2d70",
   898 => x"882a7188",
   899 => x"2b077083",
   900 => x"ffff0683",
   901 => x"ffe0800c",
   902 => x"5252028c",
   903 => x"050d0402",
   904 => x"f8050d73",
   905 => x"70902b71",
   906 => x"902a0783",
   907 => x"ffe0800c",
   908 => x"52028805",
   909 => x"0d040000",
   910 => x"00ffffff",
   911 => x"ff00ffff",
   912 => x"ffff00ff",
   913 => x"ffffff00",
   914 => x"46415431",
   915 => x"36202020",
   916 => x"00000000",
   917 => x"46415433",
   918 => x"32202020",
   919 => x"00000000",
	others => x"00000000"
);

begin

mem_busy<=mem_readEnable; -- we're done on the cycle after we serve the read request

process (clk, areset)
begin
		if areset = '1' then
		elsif (clk'event and clk = '1') then
			if (mem_writeEnable = '1') then
				ram(to_integer(unsigned(mem_addr(maxAddrBit downto minAddrBit)))) := mem_write;
			end if;
		if (mem_readEnable = '1') then
			mem_read <= ram(to_integer(unsigned(mem_addr(maxAddrBit downto minAddrBit))));
		end if;
	end if;
end process;




end arch;

